module riscv ( clk, rst, inst_i, inst_addr_o, data_i, data_we_o, 
        data_ce_o, data_addr_o, data_o );
  input [31:0] inst_i;
  output [31:0] inst_addr_o;
  input [31:0] data_i;
  output [31:0] data_addr_o;
  output [31:0] data_o;
  input clk, rst;
  output data_ce_o, data_we_o;

  CKINVDCx10_ASAP7_75t_R U1 ( .A(rst), .Y(data_ce_o) );
   DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_0_ ( .D(IF__n155), .CLK(clk), .SETN(IF__n65), 
        .RESETN(IF__n67), .QN(IF__n257) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_31_ ( .D(IF__n36), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n230) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_1_ ( .D(IF__n96), .CLK(clk), .SETN(IF__n65), 
        .RESETN(IF__n67), .QN(IF__n256) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_2_ ( .D(IF__n6), .CLK(clk), .SETN(IF__IF__n67), 
        .RESETN(IF__IF__n65), .QN(IF__n255) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_3_ ( .D(IF__n156), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n254) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_4_ ( .D(IF__n56), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n253) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_5_ ( .D(IF__n19), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n252) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_6_ ( .D(IF__n157), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n251) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_7_ ( .D(IF__n9), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n250) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_8_ ( .D(IF__n11), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n249) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_10_ ( .D(IF__n43), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(inst_addr_o[10]) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_11_ ( .D(IF__n38), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(inst_addr_o[11]) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_12_ ( .D(IF__n33), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n247) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_13_ ( .D(IF__n44), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n246) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_14_ ( .D(IF__n37), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n245) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_15_ ( .D(IF__n41), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n244) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_16_ ( .D(IF__n160), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n243) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_17_ ( .D(IF__n49), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n242) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_18_ ( .D(IF__n35), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n241) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_19_ ( .D(IF__n42), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n240) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_20_ ( .D(IF__n34), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n239) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_21_ ( .D(IF__n32), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n238) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_22_ ( .D(IF__n20), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n237) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_23_ ( .D(IF__n48), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n236) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_24_ ( .D(IF__n40), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n235) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_25_ ( .D(IF__n8), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n234) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_26_ ( .D(IF__n15), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(inst_addr_o[26]) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_27_ ( .D(IF__n91), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(inst_addr_o[27]) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_28_ ( .D(IF__n172), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n233) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_29_ ( .D(IF__n10), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n232) );
  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_30_ ( .D(IF__n84), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n231) );
  CKINVDCx10_ASAP7_75t_R IF___U66 ( .A(rst), .Y(IF__n65) );
 // IF_DW01_add_2 IF___add_17 ( .A({inst_addr_o[31:26], n28, inst_addr_o[24:23], n237, n151, 
 //       n150, n201, inst_addr_o[18], n193, n178, inst_addr_o[15:14], n246, n109, 
 //       inst_addr_o[11:10], n248, n30, n250, n251, n252, n253, n45, inst_addr_o[2], 
 //       n141, n137}), .SUM(seq_addr) );
  BUFx2_ASAP7_75t_R IF_DW01___U0 ( .A(inst_addr_o[31]), .Y(seq_addr[31]) );
  BUFx2_ASAP7_75t_R IF_DW01___U1 ( .A(inst_addr_o[30]), .Y(seq_addr[30]) );
  BUFx2_ASAP7_75t_R IF_DW01___U2 ( .A(inst_addr_o[29]), .Y(seq_addr[29]) );
  BUFx2_ASAP7_75t_R IF_DW01___U3 ( .A(inst_addr_o[28]), .Y(seq_addr[28]) );
  BUFx2_ASAP7_75t_R IF_DW01___U4 ( .A(inst_addr_o[27]), .Y(seq_addr[27]) );
  BUFx2_ASAP7_75t_R IF_DW01___U5 ( .A(inst_addr_o[26]), .Y(seq_addr[26]) );
  BUFx2_ASAP7_75t_R IF_DW01___U6 ( .A(IF__n28), .Y(seq_addr[25]) );
  BUFx2_ASAP7_75t_R IF_DW01___U7 ( .A(inst_addr_o[24]), .Y(seq_addr[24]) );
  BUFx2_ASAP7_75t_R IF_DW01___U8 ( .A(inst_addr_o[23]), .Y(seq_addr[23]) );
  BUFx2_ASAP7_75t_R IF_DW01___U9 ( .A(IF__n237), .Y(seq_addr[22]) );
  BUFx2_ASAP7_75t_R IF_DW01___U10 ( .A(IF__n151), .Y(seq_addr[21]) );
  BUFx2_ASAP7_75t_R IF_DW01___U11 ( .A(IF__n150), .Y(seq_addr[20]) );
  BUFx2_ASAP7_75t_R IF_DW01___U12 ( .A(IF__n201), .Y(seq_addr[19]) );
  BUFx2_ASAP7_75t_R IF_DW01___U13 ( .A(inst_addr_o[18]), .Y(seq_addr[18]) );
  BUFx2_ASAP7_75t_R IF_DW01___U14 ( .A(IF__n193), .Y(seq_addr[17]) );
  BUFx2_ASAP7_75t_R IF_DW01___U15 ( .A(IF__n178), .Y(seq_addr[16]) );
  BUFx2_ASAP7_75t_R IF_DW01___U16 ( .A(inst_addr_o[15]), .Y(seq_addr[15]) );
  BUFx2_ASAP7_75t_R IF_DW01___U17 ( .A(inst_addr_o[14]), .Y(seq_addr[14]) );
  BUFx2_ASAP7_75t_R IF_DW01___U18 ( .A(IF__n246), .Y(seq_addr[13]) );
  BUFx2_ASAP7_75t_R IF_DW01___U19 ( .A(IF__n109), .Y(seq_addr[12]) );
  BUFx2_ASAP7_75t_R IF_DW01___U20 ( .A(inst_addr_o[11]), .Y(seq_addr[11]) );
  BUFx2_ASAP7_75t_R IF_DW01___U21 ( .A(inst_addr_o[10]), .Y(seq_addr[10]) );
  BUFx2_ASAP7_75t_R IF_DW01___U22 ( .A(IF__n248), .Y(seq_addr[9]) );
  BUFx2_ASAP7_75t_R IF_DW01___U23 ( .A(IF__n30), .Y(seq_addr[8]) );
  BUFx2_ASAP7_75t_R IF_DW01___U24 ( .A(IF__n250), .Y(seq_addr[7]) );
  BUFx2_ASAP7_75t_R IF_DW01___U25 ( .A(IF__n251), .Y(seq_addr[6]) );
  BUFx2_ASAP7_75t_R IF_DW01___U26 ( .A(IF__n252), .Y(seq_addr[5]) );
  BUFx2_ASAP7_75t_R IF_DW01___U27 ( .A(IF__n253), .Y(seq_addr[4]) );
  BUFx2_ASAP7_75t_R IF_DW01___U28 ( .A(IF__n45), .Y(seq_addr[3]) );
  BUFx2_ASAP7_75t_R IF_DW01___U29 ( .A(inst_addr_o[2]), .Y(seq_addr[2]) );
  BUFx2_ASAP7_75t_R IF_DW01___U30 ( .A(IF__n141), .Y(seq_addr[1]) );
  BUFx2_ASAP7_75t_R IF_DW01___U31 ( .A(IF__n137), .Y(seq_addr[0]) );

  DFFASRHQNx1_ASAP7_75t_R IF___in_addr_reg_9_ ( .D(IF__n7), .CLK(clk), .SETN(IF__n67), 
        .RESETN(IF__n65), .QN(IF__n248) );
  TIEHIx1_ASAP7_75t_R IF___U3 ( .H(IF__n67) );
  NAND2xp5_ASAP7_75t_R IF___U4 ( .A(EX_branch_addr[0]), .B(IF__n138), .Y(IF__n57) );
  NAND2xp5_ASAP7_75t_R IF___U5 ( .A(EX_branch_addr[2]), .B(IF__n138), .Y(IF__n60) );
  NOR2x1_ASAP7_75t_R IF___U6 ( .A(IF__n2), .B(IF__n3), .Y(IF__n9) );
  
  AND2x2_ASAP7_75t_R IF___U7 ( .A(IF__n100), .B(seq_addr[7]), .Y(IF__n2) );
  OR2x2_ASAP7_75t_R IF___U8 ( .A(IF__n21), .B(IF__n22), .Y(IF__n3) );
  HB1xp67_ASAP7_75t_R IF___U9 ( .A(IF__n95), .Y(IF__n4) );
  BUFx6f_ASAP7_75t_R IF___U10 ( .A(IF__n222), .Y(IF__n138) );
  AND2x2_ASAP7_75t_R IF___U11 ( .A(IF__n125), .B(IF__n124), .Y(IF__n5) );
  AND2x2_ASAP7_75t_R IF___U12 ( .A(IF__n126), .B(IF__n5), .Y(IF__n10) );
  NAND2xp5_ASAP7_75t_R IF___U13 ( .A(EX_branch_addr[6]), .B(IF__n69), .Y(IF__n101) );
  AND3x2_ASAP7_75t_R IF___U14 ( .A(IF__IF__n60), .B(IF__IF__n61), .C(IF__IF__n62), .Y(IF__n6) );
  AND3x2_ASAP7_75t_R IF___U15 ( .A(IF__n53), .B(IF__n54), .C(IF__n55), .Y(IF__n7) );
  AND2x2_ASAP7_75t_R IF___U16 ( .A(IF__n76), .B(IF__n23), .Y(IF__n8) );
  NOR3xp33_ASAP7_75t_R IF___U17 ( .A(IF__n12), .B(IF__n13), .C(IF__n14), .Y(IF__n11) );
  AND2x2_ASAP7_75t_R IF___U18 ( .A(EX_branch_addr[8]), .B(IF__n69), .Y(IF__n12) );
  AND2x2_ASAP7_75t_R IF___U19 ( .A(IF__n144), .B(inst_addr_o[8]), .Y(IF__n13) );
  AND2x2_ASAP7_75t_R IF___U20 ( .A(seq_addr[8]), .B(IF__n100), .Y(IF__n14) );
  NAND2xp5_ASAP7_75t_R IF___U21 ( .A(IF__n119), .B(IF__n118), .Y(IF__n79) );
  NAND2xp67_ASAP7_75t_R IF___U22 ( .A(IF__n144), .B(inst_addr_o[27]), .Y(IF__n121) );
  NAND2xp5_ASAP7_75t_R IF___U23 ( .A(IF__n121), .B(IF__n120), .Y(IF__n97) );
  NOR2xp67_ASAP7_75t_R IF___U24 ( .A(IF__n85), .B(IF__n90), .Y(IF__n84) );
  NOR3xp33_ASAP7_75t_R IF___U25 ( .A(IF__n16), .B(IF__n17), .C(IF__n18), .Y(IF__n15) );
  AND2x2_ASAP7_75t_R IF___U26 ( .A(IF__n69), .B(EX_branch_addr[26]), .Y(IF__n16) );
  AND2x2_ASAP7_75t_R IF___U27 ( .A(IF__n100), .B(seq_addr[26]), .Y(IF__n17) );
  AND2x2_ASAP7_75t_R IF___U28 ( .A(IF__n144), .B(inst_addr_o[26]), .Y(IF__n18) );
  AND3x1_ASAP7_75t_R IF___U29 ( .A(IF__n4), .B(IF__n94), .C(IF__n93), .Y(IF__n19) );
  NAND2xp5_ASAP7_75t_R IF___U30 ( .A(IF__n144), .B(inst_addr_o[5]), .Y(IF__n94) );
  NAND2xp5_ASAP7_75t_R IF___U31 ( .A(EX_branch_addr[5]), .B(IF__n69), .Y(IF__n93) );
  AND3x1_ASAP7_75t_R IF___U32 ( .A(IF__n127), .B(IF__n128), .C(IF__n129), .Y(IF__n20) );
  NAND2xp5_ASAP7_75t_R IF___U33 ( .A(IF__n144), .B(IF__n180), .Y(IF__n128) );
  AND2x2_ASAP7_75t_R IF___U34 ( .A(IF__n144), .B(IF__n83), .Y(IF__n21) );
  AND2x2_ASAP7_75t_R IF___U35 ( .A(EX_branch_addr[7]), .B(IF__n69), .Y(IF__n22) );
  NAND2xp33_ASAP7_75t_R IF___U36 ( .A(seq_addr[29]), .B(IF__n100), .Y(IF__n126) );
  NAND2xp5_ASAP7_75t_R IF___U37 ( .A(IF__n144), .B(inst_addr_o[29]), .Y(IF__n125) );
  NAND2xp5_ASAP7_75t_R IF___U38 ( .A(IF__n137), .B(IF__n144), .Y(IF__n58) );
  AND2x2_ASAP7_75t_R IF___U39 ( .A(IF__n75), .B(IF__n74), .Y(IF__n23) );
  AND2x6_ASAP7_75t_R IF___U40 ( .A(IF__n24), .B(IF__n133), .Y(IF__n222) );
  AND2x2_ASAP7_75t_R IF___U41 ( .A(EX_PCSrc), .B(IF__n25), .Y(IF__n24) );
  INVx1_ASAP7_75t_R IF___U42 ( .A(IF__n134), .Y(IF__n25) );
  BUFx16f_ASAP7_75t_R IF___U43 ( .A(IF__n222), .Y(IF__n69) );
  CKINVDCx16_ASAP7_75t_R IF___U44 ( .A(IF__n99), .Y(IF__n100) );
  CKINVDCx10_ASAP7_75t_R IF___U45 ( .A(IF__n158), .Y(IF__n99) );
  AND2x6_ASAP7_75t_R IF___U46 ( .A(IF__n175), .B(IF__n51), .Y(IF__n158) );
  HB1xp67_ASAP7_75t_R IF___U47 ( .A(IF__n234), .Y(IF__n26) );
  BUFx2_ASAP7_75t_R IF___U48 ( .A(IF__n234), .Y(IF__n27) );
  BUFx6f_ASAP7_75t_R IF___U49 ( .A(IF__n234), .Y(IF__n28) );
  HB1xp67_ASAP7_75t_R IF___U50 ( .A(IF__n234), .Y(inst_addr_o[25]) );
  BUFx6f_ASAP7_75t_R IF___U51 ( .A(IF__n249), .Y(IF__n30) );
  BUFx4f_ASAP7_75t_R IF___U52 ( .A(IF__n249), .Y(inst_addr_o[8]) );
  AO222x2_ASAP7_75t_R IF___U53 ( .A1(IF__n69), .A2(EX_branch_addr[21]), .B1(IF__n144), .B2(
        n154), .C1(seq_addr[21]), .C2(IF__n100), .Y(IF__n115) );
  INVx1_ASAP7_75t_R IF___U54 ( .A(IF__n115), .Y(IF__n32) );
  AO222x2_ASAP7_75t_R IF___U55 ( .A1(IF__n69), .A2(EX_branch_addr[12]), .B1(IF__n144), .B2(
        n110), .C1(seq_addr[12]), .C2(IF__n100), .Y(IF__n71) );
  INVx1_ASAP7_75t_R IF___U56 ( .A(IF__n71), .Y(IF__n33) );
  AO222x2_ASAP7_75t_R IF___U57 ( .A1(IF__n69), .A2(EX_branch_addr[20]), .B1(IF__n144), .B2(
        inst_addr_o[20]), .C1(seq_addr[20]), .C2(IF__n100), .Y(IF__n82) );
  INVx1_ASAP7_75t_R IF___U58 ( .A(IF__n82), .Y(IF__n34) );
  AO222x2_ASAP7_75t_R IF___U59 ( .A1(IF__n69), .A2(EX_branch_addr[18]), .B1(IF__n144), .B2(
        inst_addr_o[18]), .C1(seq_addr[18]), .C2(IF__n100), .Y(IF__n87) );
  INVx1_ASAP7_75t_R IF___U60 ( .A(IF__n87), .Y(IF__n35) );
  AO222x2_ASAP7_75t_R IF___U61 ( .A1(IF__n69), .A2(EX_branch_addr[31]), .B1(IF__n100), .B2(
        seq_addr[31]), .C1(IF__n144), .C2(inst_addr_o[31]), .Y(IF__n112) );
  INVx1_ASAP7_75t_R IF___U62 ( .A(IF__n112), .Y(IF__n36) );
  AO222x2_ASAP7_75t_R IF___U63 ( .A1(IF__n69), .A2(EX_branch_addr[14]), .B1(IF__n144), .B2(
        inst_addr_o[14]), .C1(seq_addr[14]), .C2(IF__n100), .Y(IF__n80) );
  INVx1_ASAP7_75t_R IF___U64 ( .A(IF__n80), .Y(IF__n37) );
  AO222x2_ASAP7_75t_R IF___U65 ( .A1(IF__n69), .A2(EX_branch_addr[11]), .B1(IF__n144), .B2(
        inst_addr_o[11]), .C1(seq_addr[11]), .C2(IF__n100), .Y(IF__n117) );
  INVx1_ASAP7_75t_R IF___U67 ( .A(IF__n117), .Y(IF__n38) );
  BUFx12f_ASAP7_75t_R IF___U68 ( .A(IF__n244), .Y(inst_addr_o[15]) );
  AO222x2_ASAP7_75t_R IF___U69 ( .A1(IF__n69), .A2(EX_branch_addr[24]), .B1(IF__n144), .B2(
        inst_addr_o[24]), .C1(seq_addr[24]), .C2(IF__n100), .Y(IF__n114) );
  INVx1_ASAP7_75t_R IF___U70 ( .A(IF__n114), .Y(IF__n40) );
  AO222x2_ASAP7_75t_R IF___U71 ( .A1(IF__n69), .A2(EX_branch_addr[15]), .B1(IF__n144), .B2(
        inst_addr_o[15]), .C1(seq_addr[15]), .C2(IF__n100), .Y(IF__n88) );
  INVx1_ASAP7_75t_R IF___U72 ( .A(IF__n88), .Y(IF__n41) );
  AO222x2_ASAP7_75t_R IF___U73 ( .A1(IF__n69), .A2(EX_branch_addr[19]), .B1(IF__n144), .B2(
        inst_addr_o[19]), .C1(seq_addr[19]), .C2(IF__n100), .Y(IF__n64) );
  INVx1_ASAP7_75t_R IF___U74 ( .A(IF__n64), .Y(IF__n42) );
  AO222x2_ASAP7_75t_R IF___U75 ( .A1(IF__n69), .A2(EX_branch_addr[10]), .B1(IF__n144), .B2(IF__n66), .C1(seq_addr[10]), .C2(IF__n100), .Y(IF__n116) );
  INVx1_ASAP7_75t_R IF___U76 ( .A(IF__n116), .Y(IF__n43) );
  AO222x2_ASAP7_75t_R IF___U77 ( .A1(IF__n69), .A2(EX_branch_addr[13]), .B1(IF__n144), .B2(
        inst_addr_o[13]), .C1(seq_addr[13]), .C2(IF__n100), .Y(IF__n98) );
  INVx1_ASAP7_75t_R IF___U78 ( .A(IF__n98), .Y(IF__n44) );
  BUFx6f_ASAP7_75t_R IF___U79 ( .A(IF__n254), .Y(IF__n45) );
  BUFx2_ASAP7_75t_R IF___U80 ( .A(IF__n254), .Y(IF__n46) );
  BUFx3_ASAP7_75t_R IF___U81 ( .A(IF__n254), .Y(inst_addr_o[3]) );
  CKINVDCx12_ASAP7_75t_R IF___U82 ( .A(IF__n68), .Y(IF__n144) );
  BUFx3_ASAP7_75t_R IF___U83 ( .A(inst_addr_o[7]), .Y(IF__n83) );
  AO222x2_ASAP7_75t_R IF___U84 ( .A1(IF__n69), .A2(EX_branch_addr[23]), .B1(IF__n144), .B2(
        inst_addr_o[23]), .C1(seq_addr[23]), .C2(IF__n100), .Y(IF__n113) );
  INVx1_ASAP7_75t_R IF___U85 ( .A(IF__n113), .Y(IF__n48) );
  AO222x2_ASAP7_75t_R IF___U86 ( .A1(IF__n69), .A2(EX_branch_addr[17]), .B1(IF__n144), .B2(
        inst_addr_o[17]), .C1(seq_addr[17]), .C2(IF__n100), .Y(IF__n86) );
  INVx1_ASAP7_75t_R IF___U87 ( .A(IF__n86), .Y(IF__n49) );
  BUFx2_ASAP7_75t_R IF___U88 ( .A(IF__n242), .Y(IF__n145) );
  HB1xp67_ASAP7_75t_R IF___U89 ( .A(IF__n209), .Y(inst_addr_o[16]) );
  INVxp33_ASAP7_75t_R IF___U90 ( .A(IF__n106), .Y(IF__n108) );
  BUFx6f_ASAP7_75t_R IF___U91 ( .A(IF__n189), .Y(inst_addr_o[18]) );
  BUFx2_ASAP7_75t_R IF___U92 ( .A(IF__n241), .Y(IF__n189) );
  AND3x1_ASAP7_75t_R IF___U93 ( .A(IF__n63), .B(IF__n176), .C(IF__n177), .Y(IF__n50) );
  AND2x4_ASAP7_75t_R IF___U94 ( .A(IF__n50), .B(IF__n104), .Y(IF__n134) );
  AND2x2_ASAP7_75t_R IF___U95 ( .A(IF__n211), .B(IF__n159), .Y(IF__n51) );
  HB1xp67_ASAP7_75t_R IF___U96 ( .A(IF__n219), .Y(IF__n177) );
  INVxp33_ASAP7_75t_R IF___U97 ( .A(IF__n106), .Y(inst_addr_o[12]) );
  NAND2xp33_ASAP7_75t_R IF___U98 ( .A(IF__n100), .B(seq_addr[22]), .Y(IF__n129) );
  BUFx6f_ASAP7_75t_R IF___U99 ( .A(IF__n145), .Y(IF__n193) );
  INVxp33_ASAP7_75t_R IF___U100 ( .A(IF__n106), .Y(IF__n110) );
  INVxp67_ASAP7_75t_R IF___U101 ( .A(IF__n130), .Y(IF__n155) );
  BUFx2_ASAP7_75t_R IF___U102 ( .A(IF__n166), .Y(IF__n169) );
  BUFx2_ASAP7_75t_R IF___U103 ( .A(IF__n245), .Y(IF__n191) );
  HB1xp67_ASAP7_75t_R IF___U104 ( .A(IF__n248), .Y(inst_addr_o[9]) );
  BUFx3_ASAP7_75t_R IF___U105 ( .A(IF__n211), .Y(IF__n133) );
  NAND2xp5_ASAP7_75t_R IF___U106 ( .A(IF__n123), .B(IF__n122), .Y(IF__n90) );
  NAND2xp5_ASAP7_75t_R IF___U107 ( .A(IF__n100), .B(seq_addr[30]), .Y(IF__n123) );
  HB1xp67_ASAP7_75t_R IF___U108 ( .A(IF__n233), .Y(IF__n182) );
  BUFx3_ASAP7_75t_R IF___U109 ( .A(IF__n182), .Y(inst_addr_o[28]) );
  BUFx2_ASAP7_75t_R IF___U110 ( .A(IF__n246), .Y(inst_addr_o[13]) );
  OR2x6_ASAP7_75t_R IF___U111 ( .A(IF__n133), .B(IF__n134), .Y(IF__n68) );
  NAND2xp5_ASAP7_75t_R IF___U112 ( .A(IF__n144), .B(inst_addr_o[6]), .Y(IF__n102) );
  INVx2_ASAP7_75t_R IF___U113 ( .A(IF__n134), .Y(IF__n175) );
  NAND2xp33_ASAP7_75t_R IF___U114 ( .A(EX_branch_addr[9]), .B(IF__n69), .Y(IF__n53) );
  NAND2xp33_ASAP7_75t_R IF___U115 ( .A(IF__n144), .B(inst_addr_o[9]), .Y(IF__n54) );
  NAND2xp5_ASAP7_75t_R IF___U116 ( .A(seq_addr[9]), .B(IF__n100), .Y(IF__n55) );
  NAND2xp5_ASAP7_75t_R IF___U117 ( .A(seq_addr[6]), .B(IF__n100), .Y(IF__n103) );
  NOR2xp67_ASAP7_75t_R IF___U118 ( .A(IF__n92), .B(IF__n97), .Y(IF__n91) );
  NOR2xp67_ASAP7_75t_R IF___U119 ( .A(IF__n78), .B(IF__n79), .Y(IF__n172) );
  INVx1_ASAP7_75t_R IF___U120 ( .A(IF__n226), .Y(IF__n56) );
  HB1xp67_ASAP7_75t_R IF___U121 ( .A(IF__n250), .Y(inst_addr_o[7]) );
  NAND2xp5_ASAP7_75t_R IF___U122 ( .A(n23), .B(IF__n69), .Y(IF__n74) );
  HB1xp67_ASAP7_75t_R IF___U123 ( .A(IF__n253), .Y(inst_addr_o[4]) );
  NAND2xp5_ASAP7_75t_R IF___U124 ( .A(IF__n138), .B(EX_branch_addr[28]), .Y(IF__n118) );
  NAND2xp5_ASAP7_75t_R IF___U125 ( .A(seq_addr[0]), .B(IF__n100), .Y(IF__n59) );
  NAND3xp33_ASAP7_75t_R IF___U126 ( .A(IF__n59), .B(IF__n58), .C(IF__n57), .Y(IF__n229) );
  HB1xp67_ASAP7_75t_R IF___U127 ( .A(inst_addr_o[0]), .Y(IF__n137) );
  INVx1_ASAP7_75t_R IF___U128 ( .A(IF__n212), .Y(IF__n211) );
  NAND2xp5_ASAP7_75t_R IF___U129 ( .A(IF__n144), .B(inst_addr_o[2]), .Y(IF__n61) );
  NAND2xp33_ASAP7_75t_R IF___U130 ( .A(seq_addr[2]), .B(IF__n100), .Y(IF__n62) );
  BUFx4f_ASAP7_75t_R IF___U131 ( .A(IF__n255), .Y(inst_addr_o[2]) );
  INVx2_ASAP7_75t_R IF___U132 ( .A(IF__n106), .Y(IF__n109) );
  BUFx6f_ASAP7_75t_R IF___U133 ( .A(IF__n191), .Y(inst_addr_o[14]) );
  HB1xp67_ASAP7_75t_R IF___U134 ( .A(IF__n167), .Y(IF__n166) );
  BUFx3_ASAP7_75t_R IF___U135 ( .A(IF__n210), .Y(IF__n209) );
  BUFx6f_ASAP7_75t_R IF___U136 ( .A(IF__n209), .Y(IF__n178) );
  INVx1_ASAP7_75t_R IF___U137 ( .A(IF__n221), .Y(IF__n63) );
  INVx2_ASAP7_75t_R IF___U138 ( .A(IF__n214), .Y(IF__n174) );
  BUFx2_ASAP7_75t_R IF___U139 ( .A(IF__n243), .Y(IF__n210) );
  HB1xp67_ASAP7_75t_R IF___U140 ( .A(inst_addr_o[10]), .Y(IF__n66) );
  HB1xp67_ASAP7_75t_R IF___U141 ( .A(IF__n251), .Y(inst_addr_o[6]) );
  BUFx6f_ASAP7_75t_R IF___U142 ( .A(IF__n208), .Y(IF__n207) );
  BUFx2_ASAP7_75t_R IF___U143 ( .A(IF__n239), .Y(IF__n148) );
  BUFx6f_ASAP7_75t_R IF___U144 ( .A(IF__n148), .Y(IF__n208) );
  NOR2xp67_ASAP7_75t_R IF___U145 ( .A(IF__n173), .B(IF__n171), .Y(IF__n72) );
  NOR3x1_ASAP7_75t_R IF___U146 ( .A(IF__n73), .B(IF__n168), .C(IF__n170), .Y(IF__n104) );
  INVx1_ASAP7_75t_R IF___U147 ( .A(IF__n72), .Y(IF__n73) );
  INVx2_ASAP7_75t_R IF___U148 ( .A(IF__n169), .Y(IF__n168) );
  INVx1_ASAP7_75t_R IF___U149 ( .A(IF__n164), .Y(IF__n171) );
  NAND2xp33_ASAP7_75t_R IF___U150 ( .A(IF__n26), .B(IF__n144), .Y(IF__n75) );
  NAND2xp33_ASAP7_75t_R IF___U151 ( .A(seq_addr[25]), .B(IF__n100), .Y(IF__n76) );
  HB1xp67_ASAP7_75t_R IF___U152 ( .A(IF__n229), .Y(IF__n130) );
  AND2x2_ASAP7_75t_R IF___U153 ( .A(IF__n144), .B(inst_addr_o[28]), .Y(IF__n78) );
  HB1xp67_ASAP7_75t_R IF___U154 ( .A(IF__n252), .Y(inst_addr_o[5]) );
  AND2x2_ASAP7_75t_R IF___U155 ( .A(IF__n69), .B(EX_branch_addr[30]), .Y(IF__n85) );
  NAND2xp33_ASAP7_75t_R IF___U156 ( .A(IF__n144), .B(inst_addr_o[30]), .Y(IF__n122) );
  AND2x2_ASAP7_75t_R IF___U157 ( .A(IF__n100), .B(seq_addr[27]), .Y(IF__n92) );
  NAND2xp33_ASAP7_75t_R IF___U158 ( .A(seq_addr[5]), .B(IF__n100), .Y(IF__n95) );
  INVx1_ASAP7_75t_R IF___U159 ( .A(IF__n228), .Y(IF__n96) );
  HB1xp67_ASAP7_75t_R IF___U160 ( .A(IF__n256), .Y(IF__n139) );
  NAND2xp5_ASAP7_75t_R IF___U161 ( .A(IF__n69), .B(EX_branch_addr[27]), .Y(IF__n120) );
  AND4x1_ASAP7_75t_R IF___U162 ( .A(inst_addr_o[5]), .B(inst_addr_o[6]), .C(inst_addr_o[7]), 
        .D(inst_addr_o[8]), .Y(IF__n216) );
  BUFx2_ASAP7_75t_R IF___U163 ( .A(IF__n230), .Y(IF__n183) );
  BUFx6f_ASAP7_75t_R IF___U164 ( .A(IF__n183), .Y(IF__n200) );
  HB1xp67_ASAP7_75t_R IF___U165 ( .A(IF__n256), .Y(inst_addr_o[1]) );
  HB1xp67_ASAP7_75t_R IF___U166 ( .A(IF__n256), .Y(IF__n142) );
  HB1xp67_ASAP7_75t_R IF___U167 ( .A(IF__n256), .Y(IF__n141) );
  INVx2_ASAP7_75t_R IF___U168 ( .A(IF__n163), .Y(IF__n170) );
  NAND3xp33_ASAP7_75t_R IF___U169 ( .A(IF__n101), .B(IF__n103), .C(IF__n102), .Y(IF__n225) );
  INVxp67_ASAP7_75t_R IF___U170 ( .A(IF__n213), .Y(IF__n105) );
  AND2x4_ASAP7_75t_R IF___U171 ( .A(inst_addr_o[30]), .B(inst_addr_o[29]), .Y(IF__n214) );
  HB1xp67_ASAP7_75t_R IF___U172 ( .A(IF__n237), .Y(IF__n180) );
  HB1xp67_ASAP7_75t_R IF___U173 ( .A(IF__n237), .Y(inst_addr_o[22]) );
  INVx2_ASAP7_75t_R IF___U174 ( .A(IF__n247), .Y(IF__n106) );
  BUFx2_ASAP7_75t_R IF___U175 ( .A(IF__n232), .Y(IF__n187) );
  HB1xp67_ASAP7_75t_R IF___U176 ( .A(stall), .Y(IF__n212) );
  BUFx6f_ASAP7_75t_R IF___U177 ( .A(IF__n187), .Y(inst_addr_o[29]) );
  BUFx6f_ASAP7_75t_R IF___U178 ( .A(IF__n196), .Y(inst_addr_o[30]) );
  INVxp67_ASAP7_75t_R IF___U179 ( .A(IF__n131), .Y(IF__n157) );
  BUFx3_ASAP7_75t_R IF___U180 ( .A(IF__n231), .Y(IF__n196) );
  HB1xp67_ASAP7_75t_R IF___U181 ( .A(IF__n218), .Y(IF__n167) );
  BUFx2_ASAP7_75t_R IF___U182 ( .A(IF__n215), .Y(IF__n163) );
  HB1xp67_ASAP7_75t_R IF___U183 ( .A(IF__n132), .Y(IF__n131) );
  HB1xp67_ASAP7_75t_R IF___U184 ( .A(IF__n225), .Y(IF__n132) );
  NAND2xp5_ASAP7_75t_R IF___U185 ( .A(IF__n100), .B(seq_addr[28]), .Y(IF__n119) );
  NAND2xp5_ASAP7_75t_R IF___U186 ( .A(IF__n138), .B(EX_branch_addr[29]), .Y(IF__n124) );
  NAND2xp5_ASAP7_75t_R IF___U187 ( .A(IF__n69), .B(EX_branch_addr[22]), .Y(IF__n127) );
  BUFx2_ASAP7_75t_R IF___U188 ( .A(IF__n197), .Y(IF__n152) );
  BUFx3_ASAP7_75t_R IF___U189 ( .A(IF__n136), .Y(IF__n135) );
  BUFx2_ASAP7_75t_R IF___U190 ( .A(IF__n257), .Y(IF__n136) );
  BUFx6f_ASAP7_75t_R IF___U191 ( .A(IF__n193), .Y(inst_addr_o[17]) );
  BUFx12f_ASAP7_75t_R IF___U192 ( .A(IF__n240), .Y(IF__n146) );
  BUFx4f_ASAP7_75t_R IF___U193 ( .A(IF__n201), .Y(inst_addr_o[19]) );
  BUFx6f_ASAP7_75t_R IF___U194 ( .A(IF__n208), .Y(inst_addr_o[20]) );
  BUFx12f_ASAP7_75t_R IF___U195 ( .A(IF__n207), .Y(IF__n150) );
  BUFx12f_ASAP7_75t_R IF___U196 ( .A(IF__n197), .Y(IF__n151) );
  BUFx2_ASAP7_75t_R IF___U197 ( .A(IF__n197), .Y(inst_addr_o[21]) );
  BUFx2_ASAP7_75t_R IF___U198 ( .A(IF__n197), .Y(IF__n154) );
  AO222x2_ASAP7_75t_R IF___U199 ( .A1(EX_branch_addr[1]), .A2(IF__n69), .B1(IF__n142), .B2(
        n144), .C1(seq_addr[1]), .C2(IF__n100), .Y(IF__n228) );
  AO222x2_ASAP7_75t_R IF___U200 ( .A1(IF__n69), .A2(EX_branch_addr[3]), .B1(IF__n144), .B2(IF__n46), .C1(seq_addr[3]), .C2(IF__n100), .Y(IF__n227) );
  INVx1_ASAP7_75t_R IF___U201 ( .A(IF__n227), .Y(IF__n156) );
  AO222x2_ASAP7_75t_R IF___U202 ( .A1(EX_branch_addr[4]), .A2(IF__n138), .B1(IF__n144), .B2(
        inst_addr_o[4]), .C1(seq_addr[4]), .C2(IF__n100), .Y(IF__n226) );
  BUFx2_ASAP7_75t_R IF___U203 ( .A(IF__n223), .Y(IF__n159) );
  AO222x2_ASAP7_75t_R IF___U204 ( .A1(EX_branch_addr[16]), .A2(IF__n69), .B1(IF__n144), .B2(
        inst_addr_o[16]), .C1(seq_addr[16]), .C2(IF__n100), .Y(IF__n224) );
  INVx1_ASAP7_75t_R IF___U205 ( .A(IF__n224), .Y(IF__n160) );
  AND4x1_ASAP7_75t_R IF___U206 ( .A(IF__n27), .B(inst_addr_o[26]), .C(inst_addr_o[27]), .D(
        inst_addr_o[28]), .Y(IF__n213) );
  BUFx3_ASAP7_75t_R IF___U207 ( .A(IF__n162), .Y(IF__n161) );
  BUFx2_ASAP7_75t_R IF___U208 ( .A(IF__n217), .Y(IF__n162) );
  AND4x1_ASAP7_75t_R IF___U209 ( .A(inst_addr_o[9]), .B(inst_addr_o[10]), .C(inst_addr_o[11]), .D(IF__n108), .Y(IF__n217) );
  AND4x1_ASAP7_75t_R IF___U210 ( .A(inst_addr_o[31]), .B(inst_addr_o[2]), .C(inst_addr_o[3]), 
        .D(inst_addr_o[4]), .Y(IF__n215) );
  BUFx3_ASAP7_75t_R IF___U211 ( .A(IF__n165), .Y(IF__n164) );
  BUFx2_ASAP7_75t_R IF___U212 ( .A(IF__n216), .Y(IF__n165) );
  AND4x1_ASAP7_75t_R IF___U213 ( .A(inst_addr_o[13]), .B(inst_addr_o[14]), .C(
        inst_addr_o[15]), .D(IF__n210), .Y(IF__n218) );
  INVx1_ASAP7_75t_R IF___U214 ( .A(IF__n161), .Y(IF__n173) );
  OR4x1_ASAP7_75t_R IF___U215 ( .A(IF__n174), .B(IF__n139), .C(IF__n105), .D(inst_addr_o[0]), .Y(
        n221) );
  BUFx2_ASAP7_75t_R IF___U216 ( .A(IF__n220), .Y(IF__n176) );
  AND4x1_ASAP7_75t_R IF___U217 ( .A(inst_addr_o[17]), .B(inst_addr_o[18]), .C(IF__n201), .D(
        inst_addr_o[20]), .Y(IF__n220) );
  AND4x1_ASAP7_75t_R IF___U218 ( .A(IF__n152), .B(inst_addr_o[22]), .C(inst_addr_o[23]), .D(
        inst_addr_o[24]), .Y(IF__n219) );
  BUFx12f_ASAP7_75t_R IF___U219 ( .A(IF__n185), .Y(inst_addr_o[23]) );
  BUFx12f_ASAP7_75t_R IF___U220 ( .A(IF__n236), .Y(IF__n185) );
  BUFx12f_ASAP7_75t_R IF___U221 ( .A(IF__n198), .Y(IF__n197) );
  BUFx12f_ASAP7_75t_R IF___U222 ( .A(IF__n238), .Y(IF__n198) );
  BUFx12f_ASAP7_75t_R IF___U223 ( .A(IF__n200), .Y(inst_addr_o[31]) );
  BUFx12f_ASAP7_75t_R IF___U224 ( .A(IF__n202), .Y(IF__n201) );
  BUFx12f_ASAP7_75t_R IF___U225 ( .A(IF__n146), .Y(IF__n202) );
  BUFx12f_ASAP7_75t_R IF___U226 ( .A(IF__n204), .Y(inst_addr_o[24]) );
  BUFx12f_ASAP7_75t_R IF___U227 ( .A(IF__n235), .Y(IF__n204) );
  BUFx6f_ASAP7_75t_R IF___U228 ( .A(IF__n206), .Y(inst_addr_o[0]) );
  BUFx4f_ASAP7_75t_R IF___U229 ( .A(IF__n135), .Y(IF__n206) );
  TIELOx1_ASAP7_75t_R IF___U230 ( .L(IF__n1) );
  INVx1_ASAP7_75t_R IF___U231 ( .A(EX_PCSrc), .Y(IF__n223) );
 DFFASRHQNx1_ASAP7_75t_R IF_ID___rs2_reg_4_ ( .D(IF_ID__n244), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n686) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rs2_reg_3_ ( .D(IF_ID__n269), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID_rs2[3]) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rs2_reg_2_ ( .D(IF_ID__n172), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID_rs2[2]) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rs2_reg_1_ ( .D(IF_ID__n232), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID_rs2[1]) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rs2_reg_0_ ( .D(IF_ID__n595), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID_rs2[0]) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_31_ ( .D(IF_ID__n158), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n687) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_30_ ( .D(IF_ID__n5), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n688) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_29_ ( .D(IF_ID__n48), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n689) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_28_ ( .D(IF_ID__n323), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n690) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_27_ ( .D(IF_ID__n181), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n691) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_26_ ( .D(IF_ID__n159), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n692) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_25_ ( .D(IF_ID__n208), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n693) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_24_ ( .D(IF_ID__n180), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n694) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_23_ ( .D(IF_ID__n7), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__IF_ID__n70), .QN(IF_ID__n695) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_22_ ( .D(IF_ID__n9), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n696) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_21_ ( .D(IF_ID__n50), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n697) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_20_ ( .D(IF_ID__n52), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n698) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_19_ ( .D(IF_ID__n46), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n699) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_18_ ( .D(IF_ID__n47), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__IF_ID__n700) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_17_ ( .D(IF_ID__n229), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__IF_ID__n701) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_16_ ( .D(IF_ID__n177), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__IF_ID__n702) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_15_ ( .D(IF_ID__n183), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__IF_ID__n703) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_14_ ( .D(IF_ID__n205), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__IF_ID__n704) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_13_ ( .D(IF_ID__n36), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__IF_ID__n705) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_12_ ( .D(IF_ID__n231), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__IF_ID__n706) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_11_ ( .D(IF_ID__n161), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__IF_ID__n707) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_10_ ( .D(IF_ID__n182), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__IF_ID__n708) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_9_ ( .D(IF_ID__n322), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__IF_ID__n709) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_8_ ( .D(IF_ID__n206), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n710) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_7_ ( .D(IF_ID__n160), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n711) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_6_ ( .D(IF_ID__n321), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n712) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_5_ ( .D(IF_ID__n207), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n713) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_4_ ( .D(IF_ID__n230), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n714) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_3_ ( .D(IF_ID__n382), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n715) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_2_ ( .D(IF_ID__n45), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n716) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_1_ ( .D(IF_ID__n44), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n717) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_addr_out_reg_0_ ( .D(IF_ID__n25), .CLK(clk), .SETN(
        n171), .RESETN(IF_ID__n70), .QN(IF_ID__n718) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_31_ ( .D(IF_ID__n26), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n719) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_30_ ( .D(IF_ID__n383), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n720) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_29_ ( .D(IF_ID__n35), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n721) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_28_ ( .D(IF_ID__n178), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n722) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_27_ ( .D(IF_ID__n33), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n723) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_26_ ( .D(IF_ID__n140), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n724) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_25_ ( .D(IF_ID__n179), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n725) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_24_ ( .D(IF_ID__n191), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n726) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_22_ ( .D(IF_ID__n233), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n728) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_21_ ( .D(IF_ID__n192), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n729) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_20_ ( .D(IF_ID__n234), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n730) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_18_ ( .D(IF_ID__n637), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n732) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_17_ ( .D(IF_ID__n638), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n733) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_16_ ( .D(IF_ID__n196), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n734) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_15_ ( .D(IF_ID__n336), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n735) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_14_ ( .D(IF_ID__n320), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n736) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_13_ ( .D(IF_ID__n34), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n737) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_12_ ( .D(IF_ID__n56), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n738) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_11_ ( .D(IF_ID__n643), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n739) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_10_ ( .D(IF_ID__n644), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n740) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_9_ ( .D(IF_ID__n645), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n741) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_8_ ( .D(IF_ID__n646), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n742) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_7_ ( .D(IF_ID__n647), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n743) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_6_ ( .D(IF_ID__n648), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n744) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_5_ ( .D(IF_ID__n433), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n745) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_4_ ( .D(IF_ID__n650), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID_inst[4]) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_3_ ( .D(IF_ID__n80), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID_inst[3]) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_2_ ( .D(IF_ID__n91), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID_inst[2]) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_1_ ( .D(IF_ID__n99), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n746) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_0_ ( .D(IF_ID__n117), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n747) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___opcode_reg_6_ ( .D(IF_ID__n655), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n672) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___opcode_reg_5_ ( .D(IF_ID__n656), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n673) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___opcode_reg_4_ ( .D(IF_ID__n657), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n674) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___opcode_reg_3_ ( .D(IF_ID__n658), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID_opcode[3]) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___opcode_reg_2_ ( .D(IF_ID__n144), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n675) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___opcode_reg_1_ ( .D(IF_ID__n236), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n676) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___opcode_reg_0_ ( .D(IF_ID__n197), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n677) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rd_reg_4_ ( .D(IF_ID__n238), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n678) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rd_reg_3_ ( .D(IF_ID__n127), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n679) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rd_reg_2_ ( .D(IF_ID__n145), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n680) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rd_reg_1_ ( .D(IF_ID__n174), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n681) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rd_reg_0_ ( .D(IF_ID__n199), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n682) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rs1_reg_3_ ( .D(IF_ID__n240), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n684) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rs1_reg_1_ ( .D(IF_ID__n247), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID_rs1[1]) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rs1_reg_0_ ( .D(IF_ID__n37), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID_rs1[0]) );
  CKINVDCx10_ASAP7_75t_R IF_ID___U173 ( .A(rst), .Y(IF_ID__n171) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rs1_reg_2_ ( .D(IF_ID__n669), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n685) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___rs1_reg_4_ ( .D(IF_ID__n667), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n683) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_19_ ( .D(IF_ID__n636), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n731) );
  DFFASRHQNx1_ASAP7_75t_R IF_ID___inst_out_reg_23_ ( .D(IF_ID__n632), .CLK(clk), .SETN(IF_ID__n171), 
        .RESETN(IF_ID__n70), .QN(IF_ID__n727) );
  TIEHIx1_ASAP7_75t_R IF_ID___U3 ( .H(IF_ID__n70) );
  AOI21xp5_ASAP7_75t_R IF_ID___U4 ( .A1(IF_ID__n213), .A2(IF_ID_opcode[2]), .B(IF_ID__n584), .Y(IF_ID__n659) );
  BUFx6f_ASAP7_75t_R IF_ID___U5 ( .A(IF_ID__n531), .Y(IF_ID__n1) );
  HB1xp67_ASAP7_75t_R IF_ID___U6 ( .A(IF_ID__n598), .Y(IF_ID__n176) );
  INVx1_ASAP7_75t_R IF_ID___U7 ( .A(IF_ID__n516), .Y(IF_ID__n2) );
  BUFx6f_ASAP7_75t_R IF_ID___U8 ( .A(IF_ID__n14), .Y(IF_ID__n15) );
  CKINVDCx10_ASAP7_75t_R IF_ID___U9 ( .A(IF_ID__n515), .Y(IF_ID__n531) );
  CKINVDCx14_ASAP7_75t_R IF_ID___U10 ( .A(IF_ID__n114), .Y(IF_ID__n515) );
  INVx4_ASAP7_75t_R IF_ID___U11 ( .A(IF_ID__n215), .Y(IF_ID__n522) );
  AOI21xp5_ASAP7_75t_R IF_ID___U12 ( .A1(IF_ID__n516), .A2(IF_ID__n65), .B(IF_ID__n163), .Y(IF_ID__n592) );
  INVx1_ASAP7_75t_R IF_ID___U13 ( .A(IF_ID__n516), .Y(IF_ID__n528) );
  INVx1_ASAP7_75t_R IF_ID___U14 ( .A(IF_ID__n163), .Y(IF_ID__n22) );
  INVx4_ASAP7_75t_R IF_ID___U15 ( .A(IF_ID__n517), .Y(IF_ID__n532) );
  CKINVDCx6p67_ASAP7_75t_R IF_ID___U16 ( .A(IF_ID__n214), .Y(IF_ID__n521) );
  BUFx2_ASAP7_75t_R IF_ID___U17 ( .A(IF_ID__n29), .Y(IF_ID__n3) );
  BUFx3_ASAP7_75t_R IF_ID___U18 ( .A(IF_ID__n30), .Y(IF_ID__n4) );
  INVx3_ASAP7_75t_R IF_ID___U19 ( .A(IF_ID__n69), .Y(IF_ID__n29) );
  AND2x2_ASAP7_75t_R IF_ID___U20 ( .A(inst_i[21]), .B(IF_ID__n28), .Y(IF_ID__n558) );
  BUFx4f_ASAP7_75t_R IF_ID___U21 ( .A(IF_ID__n30), .Y(IF_ID__n21) );
  INVx2_ASAP7_75t_R IF_ID___U22 ( .A(IF_ID__n221), .Y(IF_ID__n402) );
  BUFx3_ASAP7_75t_R IF_ID___U23 ( .A(IF_ID__n576), .Y(IF_ID__n221) );
  CKINVDCx10_ASAP7_75t_R IF_ID___U24 ( .A(IF_ID__n112), .Y(IF_ID__n529) );
  INVx5_ASAP7_75t_R IF_ID___U25 ( .A(IF_ID__n529), .Y(IF_ID__n13) );
  INVx13_ASAP7_75t_R IF_ID___U26 ( .A(IF_ID__n12), .Y(IF_ID__n518) );
  BUFx16f_ASAP7_75t_R IF_ID___U27 ( .A(IF_ID__n114), .Y(IF_ID__n12) );
  INVx6_ASAP7_75t_R IF_ID___U28 ( .A(IF_ID__n518), .Y(IF_ID__n527) );
  AND2x2_ASAP7_75t_R IF_ID___U29 ( .A(IF_ID__n42), .B(IF_ID__n43), .Y(IF_ID__n5) );
  AO22x1_ASAP7_75t_R IF_ID___U30 ( .A1(inst_addr_o[23]), .A2(IF_ID__n21), .B1(
        IF_ID_inst_addr[23]), .B2(IF_ID__n11), .Y(IF_ID__n6) );
  CKINVDCx8_ASAP7_75t_R IF_ID___U31 ( .A(IF_ID__n69), .Y(IF_ID__n30) );
  AO22x2_ASAP7_75t_R IF_ID___U32 ( .A1(inst_addr_o[21]), .A2(IF_ID__n21), .B1(
        IF_ID_inst_addr[21]), .B2(IF_ID__n518), .Y(IF_ID__n603) );
  INVxp67_ASAP7_75t_R IF_ID___U33 ( .A(IF_ID__n6), .Y(IF_ID__n7) );
  INVx1_ASAP7_75t_R IF_ID___U34 ( .A(IF_ID__n584), .Y(IF_ID__n406) );
  AO22x2_ASAP7_75t_R IF_ID___U35 ( .A1(inst_i[28]), .A2(IF_ID__n3), .B1(IF_ID_inst[28]), .B2(
        n214), .Y(IF_ID__n627) );
  INVx1_ASAP7_75t_R IF_ID___U36 ( .A(IF_ID__n627), .Y(IF_ID__n178) );
  AO22x1_ASAP7_75t_R IF_ID___U37 ( .A1(IF_ID__n8), .A2(IF_ID__n21), .B1(IF_ID_inst[25]), .B2(IF_ID__n13), .Y(
        n630) );
  CKINVDCx20_ASAP7_75t_R IF_ID___U38 ( .A(IF_ID__n32), .Y(IF_ID__n8) );
  INVx2_ASAP7_75t_R IF_ID___U39 ( .A(IF_ID__n582), .Y(IF_ID__n407) );
  INVx2_ASAP7_75t_R IF_ID___U40 ( .A(IF_ID__n570), .Y(IF_ID__n404) );
  BUFx2_ASAP7_75t_R IF_ID___U41 ( .A(IF_ID__n153), .Y(IF_ID__n152) );
  AND2x2_ASAP7_75t_R IF_ID___U42 ( .A(IF_ID__n40), .B(IF_ID__n41), .Y(IF_ID__n9) );
  BUFx6f_ASAP7_75t_R IF_ID___U43 ( .A(IF_ID__n216), .Y(IF_ID__n10) );
  INVx4_ASAP7_75t_R IF_ID___U44 ( .A(IF_ID__n216), .Y(IF_ID__n23) );
  BUFx2_ASAP7_75t_R IF_ID___U45 ( .A(IF_ID__n76), .Y(IF_ID__n116) );
  INVx2_ASAP7_75t_R IF_ID___U46 ( .A(IF_ID__n11), .Y(IF_ID__n76) );
  HB1xp67_ASAP7_75t_R IF_ID___U47 ( .A(IF_ID__n659), .Y(IF_ID__n144) );
  AO22x2_ASAP7_75t_R IF_ID___U48 ( .A1(inst_i[27]), .A2(IF_ID__n21), .B1(IF_ID_inst[27]), .B2(
        n533), .Y(IF_ID__n628) );
  HB1xp67_ASAP7_75t_R IF_ID___U49 ( .A(IF_ID__n596), .Y(IF_ID__n79) );
  HB1xp67_ASAP7_75t_R IF_ID___U50 ( .A(IF_ID__n615), .Y(IF_ID__n134) );
  HB1xp67_ASAP7_75t_R IF_ID___U51 ( .A(IF_ID__n610), .Y(IF_ID__n110) );
  AOI22x1_ASAP7_75t_R IF_ID___U52 ( .A1(inst_i[13]), .A2(IF_ID__n15), .B1(IF_ID__n215), .B2(
        IF_ID_inst[13]), .Y(IF_ID__n34) );
  BUFx12f_ASAP7_75t_R IF_ID___U53 ( .A(IF_ID__n10), .Y(IF_ID__n115) );
  HB1xp67_ASAP7_75t_R IF_ID___U54 ( .A(IF_ID__n607), .Y(IF_ID__n147) );
  HB1xp67_ASAP7_75t_R IF_ID___U55 ( .A(IF_ID__n621), .Y(IF_ID__n89) );
  HB1xp67_ASAP7_75t_R IF_ID___U56 ( .A(IF_ID__n608), .Y(IF_ID__n102) );
  HB1xp67_ASAP7_75t_R IF_ID___U57 ( .A(IF_ID__n620), .Y(IF_ID__n149) );
  INVx6_ASAP7_75t_R IF_ID___U58 ( .A(IF_ID__n531), .Y(IF_ID__n11) );
  HB1xp67_ASAP7_75t_R IF_ID___U59 ( .A(IF_ID__n609), .Y(IF_ID__n98) );
  BUFx16f_ASAP7_75t_R IF_ID___U60 ( .A(IF_ID__n512), .Y(IF_ID__n214) );
  INVx6_ASAP7_75t_R IF_ID___U61 ( .A(IF_ID__n115), .Y(IF_ID__n512) );
  BUFx16f_ASAP7_75t_R IF_ID___U62 ( .A(IF_ID__n216), .Y(IF_ID__n114) );
  INVx2_ASAP7_75t_R IF_ID___U63 ( .A(IF_ID__n514), .Y(IF_ID__n526) );
  AO22x2_ASAP7_75t_R IF_ID___U64 ( .A1(IF_ID__n14), .A2(inst_addr_o[19]), .B1(
        IF_ID_inst_addr[19]), .B2(IF_ID__n518), .Y(IF_ID__n605) );
  INVx3_ASAP7_75t_R IF_ID___U65 ( .A(IF_ID__n164), .Y(IF_ID__n400) );
  BUFx3_ASAP7_75t_R IF_ID___U66 ( .A(IF_ID__n556), .Y(IF_ID__n165) );
  INVx2_ASAP7_75t_R IF_ID___U67 ( .A(IF_ID__n558), .Y(IF_ID__n358) );
  BUFx4f_ASAP7_75t_R IF_ID___U68 ( .A(IF_ID__n572), .Y(IF_ID__n222) );
  INVx2_ASAP7_75t_R IF_ID___U69 ( .A(IF_ID__n222), .Y(IF_ID__n403) );
  BUFx12f_ASAP7_75t_R IF_ID___U70 ( .A(IF_ID__n23), .Y(IF_ID__n112) );
  INVx2_ASAP7_75t_R IF_ID___U71 ( .A(IF_ID__n213), .Y(IF_ID__n525) );
  INVx2_ASAP7_75t_R IF_ID___U72 ( .A(IF_ID__n115), .Y(IF_ID__n513) );
  INVx1_ASAP7_75t_R IF_ID___U73 ( .A(IF_ID__n103), .Y(IF_ID__n182) );
  BUFx2_ASAP7_75t_R IF_ID___U74 ( .A(IF_ID__n104), .Y(IF_ID__n103) );
  INVx2_ASAP7_75t_R IF_ID___U75 ( .A(IF_ID__n170), .Y(IF_ID__n363) );
  AND2x4_ASAP7_75t_R IF_ID___U76 ( .A(inst_i[7]), .B(IF_ID__n29), .Y(IF_ID__n570) );
  BUFx6f_ASAP7_75t_R IF_ID___U77 ( .A(IF_ID__n49), .Y(IF_ID__n216) );
  INVx3_ASAP7_75t_R IF_ID___U78 ( .A(IF_ID__n168), .Y(IF_ID__n362) );
  BUFx3_ASAP7_75t_R IF_ID___U79 ( .A(IF_ID__n590), .Y(IF_ID__n169) );
  NOR2xp67_ASAP7_75t_R IF_ID___U80 ( .A(IF_ID__n27), .B(IF_ID__n219), .Y(IF_ID__n667) );
  BUFx3_ASAP7_75t_R IF_ID___U81 ( .A(IF_ID__n31), .Y(IF_ID__n14) );
  INVx1_ASAP7_75t_R IF_ID___U82 ( .A(IF_ID__n150), .Y(IF_ID__n206) );
  BUFx2_ASAP7_75t_R IF_ID___U83 ( .A(IF_ID__n151), .Y(IF_ID__n150) );
  INVx1_ASAP7_75t_R IF_ID___U84 ( .A(IF_ID__n94), .Y(IF_ID__n161) );
  BUFx2_ASAP7_75t_R IF_ID___U85 ( .A(IF_ID__n95), .Y(IF_ID__n94) );
  INVx1_ASAP7_75t_R IF_ID___U86 ( .A(IF_ID__n84), .Y(IF_ID__n140) );
  BUFx2_ASAP7_75t_R IF_ID___U87 ( .A(IF_ID__n85), .Y(IF_ID__n84) );
  BUFx2_ASAP7_75t_R IF_ID___U88 ( .A(IF_ID__n83), .Y(IF_ID__n82) );
  INVx3_ASAP7_75t_R IF_ID___U89 ( .A(IF_ID__n90), .Y(IF_ID__n75) );
  AND2x4_ASAP7_75t_R IF_ID___U90 ( .A(inst_i[9]), .B(IF_ID__n30), .Y(IF_ID__n574) );
  BUFx2_ASAP7_75t_R IF_ID___U91 ( .A(IF_ID__n649), .Y(IF_ID__n433) );
  INVx2_ASAP7_75t_R IF_ID___U92 ( .A(IF_ID__n69), .Y(IF_ID__n28) );
  AO22x2_ASAP7_75t_R IF_ID___U93 ( .A1(IF_ID__n4), .A2(inst_i[31]), .B1(IF_ID_inst[31]), .B2(
        n518), .Y(IF_ID__n624) );
  AND2x2_ASAP7_75t_R IF_ID___U94 ( .A(inst_i[4]), .B(IF_ID__n29), .Y(IF_ID__n587) );
  AND2x4_ASAP7_75t_R IF_ID___U95 ( .A(inst_i[1]), .B(IF_ID__n29), .Y(IF_ID__n582) );
  BUFx4f_ASAP7_75t_R IF_ID___U96 ( .A(IF_ID__n585), .Y(IF_ID__n170) );
  AND2x4_ASAP7_75t_R IF_ID___U97 ( .A(inst_i[24]), .B(IF_ID__n30), .Y(IF_ID__n562) );
  AND2x4_ASAP7_75t_R IF_ID___U98 ( .A(inst_i[0]), .B(IF_ID__n30), .Y(IF_ID__n580) );
  BUFx3_ASAP7_75t_R IF_ID___U99 ( .A(stall), .Y(IF_ID__n534) );
  NAND2xp5_ASAP7_75t_R IF_ID___U100 ( .A(inst_addr_o[30]), .B(IF_ID__n15), .Y(IF_ID__n42) );
  AO22x2_ASAP7_75t_R IF_ID___U101 ( .A1(inst_i[29]), .A2(IF_ID__n15), .B1(IF_ID__n533), .B2(
        IF_ID_inst[29]), .Y(IF_ID__n626) );
  AND2x4_ASAP7_75t_R IF_ID___U102 ( .A(inst_i[18]), .B(IF_ID__n31), .Y(IF_ID__n568) );
  BUFx2_ASAP7_75t_R IF_ID___U103 ( .A(IF_ID__n668), .Y(IF_ID__n240) );
  CKINVDCx12_ASAP7_75t_R IF_ID___U104 ( .A(IF_ID__n124), .Y(IF_ID__n241) );
  BUFx16f_ASAP7_75t_R IF_ID___U105 ( .A(IF_ID__n203), .Y(IF_ID__n124) );
  CKINVDCx10_ASAP7_75t_R IF_ID___U106 ( .A(IF_ID__n241), .Y(IF_ID_rs1[3]) );
  BUFx2_ASAP7_75t_R IF_ID___U107 ( .A(IF_ID__n241), .Y(IF_ID__n16) );
  BUFx6f_ASAP7_75t_R IF_ID___U108 ( .A(IF_ID__n125), .Y(IF_ID__n203) );
  BUFx4f_ASAP7_75t_R IF_ID___U109 ( .A(IF_ID__n204), .Y(IF_ID__n125) );
  BUFx2_ASAP7_75t_R IF_ID___U110 ( .A(IF_ID__n55), .Y(IF_ID__n204) );
  BUFx8_ASAP7_75t_R IF_ID___U111 ( .A(IF_ID__n683), .Y(IF_ID_rs1[4]) );
  HB1xp67_ASAP7_75t_R IF_ID___U112 ( .A(IF_ID_rs1[0]), .Y(IF_ID__n19) );
  BUFx3_ASAP7_75t_R IF_ID___U113 ( .A(IF_ID__n745), .Y(IF_ID__n375) );
  HB1xp67_ASAP7_75t_R IF_ID___U114 ( .A(IF_ID_inst[3]), .Y(IF_ID__n20) );
  AND2x2_ASAP7_75t_R IF_ID___U115 ( .A(inst_i[20]), .B(IF_ID__n30), .Y(IF_ID__n556) );
  BUFx3_ASAP7_75t_R IF_ID___U116 ( .A(IF_ID__n560), .Y(IF_ID__n187) );
  BUFx2_ASAP7_75t_R IF_ID___U117 ( .A(IF_ID__n298), .Y(IF_ID__n139) );
  BUFx2_ASAP7_75t_R IF_ID___U118 ( .A(IF_ID__n299), .Y(IF_ID__n298) );
  BUFx3_ASAP7_75t_R IF_ID___U119 ( .A(IF_ID__n298), .Y(IF_ID_inst[1]) );
  NOR2xp67_ASAP7_75t_R IF_ID___U120 ( .A(IF_ID__n116), .B(IF_ID__n246), .Y(IF_ID__n27) );
  BUFx4f_ASAP7_75t_R IF_ID___U121 ( .A(IF_ID__n686), .Y(IF_ID_rs2[4]) );
  INVxp33_ASAP7_75t_R IF_ID___U122 ( .A(IF_ID__n375), .Y(IF_ID__n126) );
  AND2x2_ASAP7_75t_R IF_ID___U123 ( .A(inst_i[5]), .B(IF_ID__n30), .Y(IF_ID__n588) );
  HB1xp67_ASAP7_75t_R IF_ID___U124 ( .A(IF_ID_rs1[2]), .Y(IF_ID__n24) );
  HB1xp67_ASAP7_75t_R IF_ID___U125 ( .A(IF_ID__n136), .Y(IF_ID__n299) );
  NOR2x2_ASAP7_75t_R IF_ID___U126 ( .A(IF_flush), .B(IF_ID__n112), .Y(IF_ID__n31) );
  AND2x2_ASAP7_75t_R IF_ID___U127 ( .A(inst_i[6]), .B(IF_ID__n29), .Y(IF_ID__n590) );
  INVxp67_ASAP7_75t_R IF_ID___U128 ( .A(IF_ID__n131), .Y(IF_ID__n208) );
  INVx1_ASAP7_75t_R IF_ID___U129 ( .A(IF_ID__n623), .Y(IF_ID__n25) );
  HB1xp67_ASAP7_75t_R IF_ID___U130 ( .A(IF_ID__n132), .Y(IF_ID__n131) );
  INVx1_ASAP7_75t_R IF_ID___U131 ( .A(IF_ID__n624), .Y(IF_ID__n26) );
  HB1xp67_ASAP7_75t_R IF_ID___U132 ( .A(IF_ID__n137), .Y(IF_ID__n136) );
  NAND2xp5_ASAP7_75t_R IF_ID___U133 ( .A(IF_ID_inst_addr[22]), .B(IF_ID__n11), .Y(IF_ID__n41) );
  INVx1_ASAP7_75t_R IF_ID___U134 ( .A(IF_ID__n432), .Y(IF_ID__n246) );
  INVx2_ASAP7_75t_R IF_ID___U135 ( .A(IF_ID__n219), .Y(IF_ID__n327) );
  HB1xp67_ASAP7_75t_R IF_ID___U136 ( .A(IF_ID__n511), .Y(IF_ID__n157) );
  AND2x2_ASAP7_75t_R IF_ID___U137 ( .A(inst_i[17]), .B(IF_ID__n29), .Y(IF_ID__n566) );
  AND2x2_ASAP7_75t_R IF_ID___U138 ( .A(inst_i[23]), .B(IF_ID__n29), .Y(IF_ID__n561) );
  AND2x2_ASAP7_75t_R IF_ID___U139 ( .A(inst_i[10]), .B(IF_ID__n29), .Y(IF_ID__n576) );
  BUFx3_ASAP7_75t_R IF_ID___U140 ( .A(IF_ID__n675), .Y(IF_ID_opcode[2]) );
  HB1xp67_ASAP7_75t_R IF_ID___U141 ( .A(IF_ID__n746), .Y(IF_ID__n137) );
  BUFx2_ASAP7_75t_R IF_ID___U142 ( .A(IF_ID__n744), .Y(IF_ID__n135) );
  BUFx6f_ASAP7_75t_R IF_ID___U143 ( .A(IF_ID__n135), .Y(IF_ID__n511) );
  INVx1_ASAP7_75t_R IF_ID___U144 ( .A(stall), .Y(IF_ID__n49) );
  BUFx12f_ASAP7_75t_R IF_ID___U145 ( .A(IF_ID__n11), .Y(IF_ID__n213) );
  INVx2_ASAP7_75t_R IF_ID___U146 ( .A(IF_ID__n213), .Y(IF_ID__n524) );
  HB1xp67_ASAP7_75t_R IF_ID___U147 ( .A(IF_ID__n601), .Y(IF_ID__n132) );
  AND2x2_ASAP7_75t_R IF_ID___U148 ( .A(inst_i[15]), .B(IF_ID__n30), .Y(IF_ID__n563) );
  OR2x6_ASAP7_75t_R IF_ID___U149 ( .A(IF_flush), .B(IF_ID__n534), .Y(IF_ID__n69) );
  HB1xp67_ASAP7_75t_R IF_ID___U150 ( .A(IF_ID__n614), .Y(IF_ID__n104) );
  INVx2_ASAP7_75t_R IF_ID___U151 ( .A(IF_ID__n213), .Y(IF_ID__n523) );
  CKINVDCx20_ASAP7_75t_R IF_ID___U152 ( .A(inst_i[25]), .Y(IF_ID__n32) );
  INVx1_ASAP7_75t_R IF_ID___U153 ( .A(IF_ID__n628), .Y(IF_ID__n33) );
  INVx1_ASAP7_75t_R IF_ID___U154 ( .A(IF_ID__n626), .Y(IF_ID__n35) );
  BUFx12f_ASAP7_75t_R IF_ID___U155 ( .A(IF_ID__n114), .Y(IF_ID__n113) );
  INVx1_ASAP7_75t_R IF_ID___U156 ( .A(IF_ID__n611), .Y(IF_ID__n36) );
  HB1xp67_ASAP7_75t_R IF_ID___U157 ( .A(IF_ID__n629), .Y(IF_ID__n85) );
  HB1xp67_ASAP7_75t_R IF_ID___U158 ( .A(IF_ID__n613), .Y(IF_ID__n95) );
  INVx1_ASAP7_75t_R IF_ID___U159 ( .A(IF_ID__n671), .Y(IF_ID__n37) );
  BUFx6f_ASAP7_75t_R IF_ID___U160 ( .A(IF_ID__n685), .Y(IF_ID_rs1[2]) );
  HB1xp67_ASAP7_75t_R IF_ID___U161 ( .A(IF_ID__n20), .Y(IF_ID__n38) );
  HB1xp67_ASAP7_75t_R IF_ID___U162 ( .A(IF_ID__n617), .Y(IF_ID__n83) );
  HB1xp67_ASAP7_75t_R IF_ID___U163 ( .A(IF_ID__n616), .Y(IF_ID__n151) );
  AO22x1_ASAP7_75t_R IF_ID___U164 ( .A1(inst_i[26]), .A2(IF_ID__n29), .B1(IF_ID_inst[26]), 
        .B2(IF_ID__n533), .Y(IF_ID__n629) );
  AND2x2_ASAP7_75t_R IF_ID___U165 ( .A(inst_i[19]), .B(IF_ID__n31), .Y(IF_ID__n569) );
  AND2x2_ASAP7_75t_R IF_ID___U166 ( .A(inst_i[22]), .B(IF_ID__n30), .Y(IF_ID__n560) );
  AND2x2_ASAP7_75t_R IF_ID___U167 ( .A(inst_i[3]), .B(IF_ID__n29), .Y(IF_ID__n585) );
  AND2x2_ASAP7_75t_R IF_ID___U168 ( .A(inst_i[2]), .B(IF_ID__n30), .Y(IF_ID__n584) );
  AND2x2_ASAP7_75t_R IF_ID___U169 ( .A(inst_i[8]), .B(IF_ID__n30), .Y(IF_ID__n572) );
  AND2x2_ASAP7_75t_R IF_ID___U170 ( .A(inst_i[11]), .B(IF_ID__n28), .Y(IF_ID__n578) );
  HB1xp67_ASAP7_75t_R IF_ID___U171 ( .A(IF_ID_rs2[0]), .Y(IF_ID__n39) );
  AO22x1_ASAP7_75t_R IF_ID___U172 ( .A1(inst_addr_o[3]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[3]), .B2(IF_ID__n512), .Y(IF_ID__n621) );
  AO22x1_ASAP7_75t_R IF_ID___U174 ( .A1(inst_addr_o[17]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[17]), .B2(IF_ID__n512), .Y(IF_ID__n607) );
  NAND2xp33_ASAP7_75t_R IF_ID___U175 ( .A(inst_addr_o[22]), .B(IF_ID__n21), .Y(IF_ID__n40) );
  BUFx3_ASAP7_75t_R IF_ID___U176 ( .A(IF_ID__n447), .Y(IF_ID_inst_addr[22]) );
  NAND2xp5_ASAP7_75t_R IF_ID___U177 ( .A(IF_ID_inst_addr[30]), .B(IF_ID__n213), .Y(IF_ID__n43) );
  INVx1_ASAP7_75t_R IF_ID___U178 ( .A(IF_ID__n622), .Y(IF_ID__n44) );
  AOI22xp33_ASAP7_75t_R IF_ID___U179 ( .A1(inst_addr_o[2]), .A2(IF_ID__n15), .B1(
        IF_ID_inst_addr[2]), .B2(IF_ID__n517), .Y(IF_ID__n45) );
  INVx1_ASAP7_75t_R IF_ID___U180 ( .A(IF_ID__n605), .Y(IF_ID__n46) );
  INVx1_ASAP7_75t_R IF_ID___U181 ( .A(IF_ID__n606), .Y(IF_ID__n47) );
  HB1xp67_ASAP7_75t_R IF_ID___U182 ( .A(IF_ID__n630), .Y(IF_ID__n108) );
  INVx1_ASAP7_75t_R IF_ID___U183 ( .A(IF_ID__n597), .Y(IF_ID__n48) );
  INVxp67_ASAP7_75t_R IF_ID___U184 ( .A(IF_ID__n92), .Y(IF_ID__n180) );
  HB1xp67_ASAP7_75t_R IF_ID___U185 ( .A(IF_ID__n625), .Y(IF_ID__n153) );
  BUFx3_ASAP7_75t_R IF_ID___U186 ( .A(IF_ID__n130), .Y(IF_ID__n129) );
  INVx1_ASAP7_75t_R IF_ID___U187 ( .A(IF_ID__n603), .Y(IF_ID__n50) );
  HB1xp67_ASAP7_75t_R IF_ID___U188 ( .A(IF_ID__n684), .Y(IF_ID__n51) );
  HB1xp67_ASAP7_75t_R IF_ID___U189 ( .A(IF_ID__n93), .Y(IF_ID__n92) );
  INVx6_ASAP7_75t_R IF_ID___U190 ( .A(IF_ID__n119), .Y(IF_ID__n517) );
  INVx1_ASAP7_75t_R IF_ID___U191 ( .A(IF_ID__n604), .Y(IF_ID__n52) );
  HB1xp67_ASAP7_75t_R IF_ID___U192 ( .A(IF_ID__n602), .Y(IF_ID__n93) );
  HB1xp67_ASAP7_75t_R IF_ID___U193 ( .A(IF_ID__n619), .Y(IF_ID__n106) );
  HB1xp67_ASAP7_75t_R IF_ID___U194 ( .A(IF_ID__n612), .Y(IF_ID__n87) );
  AO22x1_ASAP7_75t_R IF_ID___U195 ( .A1(inst_addr_o[12]), .A2(IF_ID__n30), .B1(
        IF_ID_inst_addr[12]), .B2(IF_ID__n13), .Y(IF_ID__n612) );
  AO22x1_ASAP7_75t_R IF_ID___U196 ( .A1(inst_addr_o[4]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[4]), .B2(IF_ID__n513), .Y(IF_ID__n620) );
  INVxp33_ASAP7_75t_R IF_ID___U197 ( .A(IF_ID__n239), .Y(IF_ID__n319) );
  AO22x1_ASAP7_75t_R IF_ID___U198 ( .A1(inst_addr_o[6]), .A2(IF_ID__n21), .B1(IF_ID__n252), .B2(
        n533), .Y(IF_ID__n618) );
  HB1xp67_ASAP7_75t_R IF_ID___U199 ( .A(IF_ID_rs1[1]), .Y(IF_ID__n53) );
  HB1xp67_ASAP7_75t_R IF_ID___U200 ( .A(IF_ID_rs1[4]), .Y(IF_ID__n54) );
  INVxp33_ASAP7_75t_R IF_ID___U201 ( .A(IF_ID__n54), .Y(IF_ID__n212) );
  HB1xp67_ASAP7_75t_R IF_ID___U202 ( .A(IF_ID__n51), .Y(IF_ID__n55) );
  INVxp33_ASAP7_75t_R IF_ID___U203 ( .A(IF_ID_inst[4]), .Y(IF_ID__n539) );
  INVx1_ASAP7_75t_R IF_ID___U204 ( .A(IF_ID__n642), .Y(IF_ID__n56) );
  HB1xp67_ASAP7_75t_R IF_ID___U205 ( .A(IF_ID_rs2[4]), .Y(IF_ID__n57) );
  HB1xp67_ASAP7_75t_R IF_ID___U206 ( .A(IF_ID__n57), .Y(IF_ID__n58) );
  HB1xp67_ASAP7_75t_R IF_ID___U207 ( .A(IF_ID__n53), .Y(IF_ID__n60) );
  HB1xp67_ASAP7_75t_R IF_ID___U208 ( .A(IF_ID__n60), .Y(IF_ID__n61) );
  AO22x1_ASAP7_75t_R IF_ID___U209 ( .A1(inst_addr_o[20]), .A2(IF_ID__n21), .B1(
        IF_ID_inst_addr[20]), .B2(IF_ID__n518), .Y(IF_ID__n604) );
  AO22x1_ASAP7_75t_R IF_ID___U210 ( .A1(inst_addr_o[16]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[16]), .B2(IF_ID__n512), .Y(IF_ID__n608) );
  AO22x1_ASAP7_75t_R IF_ID___U211 ( .A1(inst_addr_o[31]), .A2(IF_ID__n29), .B1(
        IF_ID_inst_addr[31]), .B2(IF_ID__n515), .Y(IF_ID__n596) );
  BUFx6f_ASAP7_75t_R IF_ID___U212 ( .A(IF_ID__n562), .Y(IF_ID__n218) );
  INVx4_ASAP7_75t_R IF_ID___U213 ( .A(IF_ID__n223), .Y(IF_ID__n405) );
  BUFx6f_ASAP7_75t_R IF_ID___U214 ( .A(IF_ID__n565), .Y(IF_ID__n167) );
  INVx4_ASAP7_75t_R IF_ID___U215 ( .A(IF_ID__n166), .Y(IF_ID__n360) );
  INVx4_ASAP7_75t_R IF_ID___U216 ( .A(IF_ID__n217), .Y(IF_ID__n356) );
  AO22x1_ASAP7_75t_R IF_ID___U217 ( .A1(IF_ID__n28), .A2(inst_addr_o[18]), .B1(
        IF_ID_inst_addr[18]), .B2(IF_ID__n518), .Y(IF_ID__n606) );
  INVxp33_ASAP7_75t_R IF_ID___U218 ( .A(IF_ID__n61), .Y(IF_ID__n248) );
  INVxp33_ASAP7_75t_R IF_ID___U219 ( .A(IF_ID__n209), .Y(IF_ID__n586) );
  HB1xp67_ASAP7_75t_R IF_ID___U220 ( .A(IF_ID_rs2[1]), .Y(IF_ID__n62) );
  HB1xp67_ASAP7_75t_R IF_ID___U221 ( .A(IF_ID_rs2[3]), .Y(IF_ID__n63) );
  HB1xp67_ASAP7_75t_R IF_ID___U222 ( .A(IF_ID__n63), .Y(IF_ID__n64) );
  HB1xp67_ASAP7_75t_R IF_ID___U223 ( .A(IF_ID__n64), .Y(IF_ID__n65) );
  AO22x1_ASAP7_75t_R IF_ID___U224 ( .A1(inst_addr_o[26]), .A2(IF_ID__n21), .B1(
        IF_ID_inst_addr[26]), .B2(IF_ID__n13), .Y(IF_ID__n600) );
  AO22x1_ASAP7_75t_R IF_ID___U225 ( .A1(inst_i[12]), .A2(IF_ID__n4), .B1(IF_ID_inst[12]), .B2(
        n214), .Y(IF_ID__n642) );
  HB1xp67_ASAP7_75t_R IF_ID___U226 ( .A(IF_ID_rs2[2]), .Y(IF_ID__n66) );
  HB1xp67_ASAP7_75t_R IF_ID___U227 ( .A(IF_ID_inst[2]), .Y(IF_ID__n67) );
  HB1xp67_ASAP7_75t_R IF_ID___U228 ( .A(IF_ID__n67), .Y(IF_ID__n68) );
  INVxp67_ASAP7_75t_R IF_ID___U229 ( .A(IF_ID__n354), .Y(IF_ID__n557) );
  HB1xp67_ASAP7_75t_R IF_ID___U230 ( .A(IF_ID__n62), .Y(IF_ID__n71) );
  HB1xp67_ASAP7_75t_R IF_ID___U231 ( .A(IF_ID__n66), .Y(IF_ID__n72) );
  INVxp33_ASAP7_75t_R IF_ID___U232 ( .A(IF_ID__n72), .Y(IF_ID__n296) );
  INVxp33_ASAP7_75t_R IF_ID___U233 ( .A(IF_ID__n212), .Y(IF_ID__n73) );
  HB1xp67_ASAP7_75t_R IF_ID___U234 ( .A(IF_ID_opcode[3]), .Y(IF_ID__n209) );
  INVxp33_ASAP7_75t_R IF_ID___U235 ( .A(IF_ID__n68), .Y(IF_ID__n537) );
  INVxp33_ASAP7_75t_R IF_ID___U236 ( .A(IF_ID__n38), .Y(IF_ID__n538) );
  HB1xp67_ASAP7_75t_R IF_ID___U237 ( .A(IF_ID__n71), .Y(IF_ID__n74) );
  BUFx4f_ASAP7_75t_R IF_ID___U238 ( .A(IF_ID__n155), .Y(IF_ID__n154) );
  INVx2_ASAP7_75t_R IF_ID___U239 ( .A(IF_ID__n154), .Y(IF_ID__n245) );
  HB1xp67_ASAP7_75t_R IF_ID___U240 ( .A(IF_ID__n58), .Y(IF_ID__n155) );
  INVxp33_ASAP7_75t_R IF_ID___U241 ( .A(IF_ID__n74), .Y(IF_ID__n559) );
  INVxp67_ASAP7_75t_R IF_ID___U242 ( .A(IF_ID__n319), .Y(IF_ID__n564) );
  HB1xp67_ASAP7_75t_R IF_ID___U243 ( .A(IF_ID__n73), .Y(IF_ID__n432) );
  HB1xp67_ASAP7_75t_R IF_ID___U244 ( .A(IF_ID__n296), .Y(IF_ID__n173) );
  AO22x1_ASAP7_75t_R IF_ID___U245 ( .A1(inst_i[14]), .A2(IF_ID__n28), .B1(IF_ID_inst[14]), 
        .B2(IF_ID__n13), .Y(IF_ID__n641) );
  INVxp33_ASAP7_75t_R IF_ID___U246 ( .A(IF_ID__n24), .Y(IF_ID__n567) );
  AO22x1_ASAP7_75t_R IF_ID___U247 ( .A1(inst_addr_o[24]), .A2(IF_ID__n29), .B1(
        IF_ID_inst_addr[24]), .B2(IF_ID__n13), .Y(IF_ID__n602) );
  BUFx6f_ASAP7_75t_R IF_ID___U248 ( .A(IF_ID__n568), .Y(IF_ID__n90) );
  HB1xp67_ASAP7_75t_R IF_ID___U249 ( .A(IF_ID__n305), .Y(IF_ID__n354) );
  HB1xp67_ASAP7_75t_R IF_ID___U250 ( .A(IF_ID__n39), .Y(IF_ID__n305) );
  INVxp33_ASAP7_75t_R IF_ID___U251 ( .A(IF_ID__n19), .Y(IF_ID__n239) );
  BUFx2_ASAP7_75t_R IF_ID___U252 ( .A(IF_ID__n600), .Y(IF_ID__n77) );
  INVx3_ASAP7_75t_R IF_ID___U253 ( .A(IF_ID__n122), .Y(IF_ID__n361) );
  AO22x1_ASAP7_75t_R IF_ID___U254 ( .A1(inst_addr_o[0]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[0]), .B2(IF_ID__n518), .Y(IF_ID__n623) );
  BUFx2_ASAP7_75t_R IF_ID___U255 ( .A(IF_ID__n79), .Y(IF_ID__n78) );
  BUFx2_ASAP7_75t_R IF_ID___U256 ( .A(IF_ID__n651), .Y(IF_ID__n80) );
  BUFx2_ASAP7_75t_R IF_ID___U257 ( .A(IF_ID__n599), .Y(IF_ID__n81) );
  AO22x1_ASAP7_75t_R IF_ID___U258 ( .A1(inst_addr_o[27]), .A2(IF_ID__n14), .B1(
        IF_ID_inst_addr[27]), .B2(IF_ID__n13), .Y(IF_ID__n599) );
  INVx6_ASAP7_75t_R IF_ID___U259 ( .A(IF_ID__n111), .Y(IF_ID__n516) );
  AO22x1_ASAP7_75t_R IF_ID___U260 ( .A1(inst_addr_o[7]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[7]), .B2(IF_ID__n514), .Y(IF_ID__n617) );
  BUFx2_ASAP7_75t_R IF_ID___U261 ( .A(IF_ID__n87), .Y(IF_ID__n86) );
  BUFx2_ASAP7_75t_R IF_ID___U262 ( .A(IF_ID__n89), .Y(IF_ID__n88) );
  BUFx2_ASAP7_75t_R IF_ID___U263 ( .A(IF_ID__n652), .Y(IF_ID__n91) );
  AO22x1_ASAP7_75t_R IF_ID___U264 ( .A1(inst_addr_o[11]), .A2(IF_ID__n30), .B1(
        IF_ID_inst_addr[11]), .B2(IF_ID__n514), .Y(IF_ID__n613) );
  BUFx2_ASAP7_75t_R IF_ID___U265 ( .A(IF_ID__n618), .Y(IF_ID__n96) );
  BUFx2_ASAP7_75t_R IF_ID___U266 ( .A(IF_ID__n98), .Y(IF_ID__n97) );
  BUFx2_ASAP7_75t_R IF_ID___U267 ( .A(IF_ID__n653), .Y(IF_ID__n99) );
  BUFx2_ASAP7_75t_R IF_ID___U268 ( .A(IF_ID__n536), .Y(IF_ID__n100) );
  BUFx2_ASAP7_75t_R IF_ID___U269 ( .A(IF_ID__n102), .Y(IF_ID__n101) );
  AO22x1_ASAP7_75t_R IF_ID___U270 ( .A1(inst_addr_o[10]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[10]), .B2(IF_ID__n514), .Y(IF_ID__n614) );
  BUFx2_ASAP7_75t_R IF_ID___U271 ( .A(IF_ID__n106), .Y(IF_ID__n105) );
  AO22x1_ASAP7_75t_R IF_ID___U272 ( .A1(inst_addr_o[5]), .A2(IF_ID__n29), .B1(
        IF_ID_inst_addr[5]), .B2(IF_ID__n214), .Y(IF_ID__n619) );
  BUFx2_ASAP7_75t_R IF_ID___U273 ( .A(IF_ID__n108), .Y(IF_ID__n107) );
  BUFx2_ASAP7_75t_R IF_ID___U274 ( .A(IF_ID__n110), .Y(IF_ID__n109) );
  BUFx12f_ASAP7_75t_R IF_ID___U275 ( .A(IF_ID__n529), .Y(IF_ID__n111) );
  BUFx2_ASAP7_75t_R IF_ID___U276 ( .A(IF_ID__n654), .Y(IF_ID__n117) );
  BUFx2_ASAP7_75t_R IF_ID___U277 ( .A(IF_ID__n535), .Y(IF_ID__n118) );
  BUFx12f_ASAP7_75t_R IF_ID___U278 ( .A(IF_ID__n521), .Y(IF_ID__n119) );
  BUFx6f_ASAP7_75t_R IF_ID___U279 ( .A(IF_ID__n250), .Y(IF_ID_inst[0]) );
  BUFx3_ASAP7_75t_R IF_ID___U280 ( .A(IF_ID__n250), .Y(IF_ID__n121) );
  BUFx6f_ASAP7_75t_R IF_ID___U281 ( .A(IF_ID__n123), .Y(IF_ID__n122) );
  BUFx4f_ASAP7_75t_R IF_ID___U282 ( .A(IF_ID__n574), .Y(IF_ID__n123) );
  BUFx2_ASAP7_75t_R IF_ID___U283 ( .A(IF_ID__n663), .Y(IF_ID__n127) );
  BUFx2_ASAP7_75t_R IF_ID___U284 ( .A(IF_ID__n577), .Y(IF_ID__n128) );
  BUFx2_ASAP7_75t_R IF_ID___U285 ( .A(IF_ID__n641), .Y(IF_ID__n130) );
  BUFx2_ASAP7_75t_R IF_ID___U286 ( .A(IF_ID__n134), .Y(IF_ID__n133) );
  BUFx2_ASAP7_75t_R IF_ID___U287 ( .A(IF_ID__n492), .Y(IF_ID__n141) );
  BUFx4f_ASAP7_75t_R IF_ID___U288 ( .A(IF_ID__n580), .Y(IF_ID__n142) );
  INVx2_ASAP7_75t_R IF_ID___U289 ( .A(IF_ID__n506), .Y(IF_ID__n143) );
  BUFx2_ASAP7_75t_R IF_ID___U290 ( .A(IF_ID__n664), .Y(IF_ID__n145) );
  BUFx2_ASAP7_75t_R IF_ID___U291 ( .A(IF_ID__n147), .Y(IF_ID__n146) );
  BUFx2_ASAP7_75t_R IF_ID___U292 ( .A(IF_ID__n149), .Y(IF_ID__n148) );
  AO22x1_ASAP7_75t_R IF_ID___U293 ( .A1(inst_addr_o[1]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[1]), .B2(IF_ID__n516), .Y(IF_ID__n622) );
  BUFx12f_ASAP7_75t_R IF_ID___U294 ( .A(IF_ID__n511), .Y(IF_ID_inst[6]) );
  INVx1_ASAP7_75t_R IF_ID___U295 ( .A(IF_ID__n78), .Y(IF_ID__n158) );
  INVx1_ASAP7_75t_R IF_ID___U296 ( .A(IF_ID__n77), .Y(IF_ID__n159) );
  INVx1_ASAP7_75t_R IF_ID___U297 ( .A(IF_ID__n82), .Y(IF_ID__n160) );
  INVx3_ASAP7_75t_R IF_ID___U298 ( .A(IF_ID__n188), .Y(IF_ID__n359) );
  INVx2_ASAP7_75t_R IF_ID___U299 ( .A(IF_ID_inst[7]), .Y(IF_ID__n541) );
  BUFx4f_ASAP7_75t_R IF_ID___U300 ( .A(IF_ID__n453), .Y(IF_ID_inst_addr[18]) );
  BUFx2_ASAP7_75t_R IF_ID___U301 ( .A(IF_ID__n519), .Y(IF_ID__n162) );
  BUFx4f_ASAP7_75t_R IF_ID___U302 ( .A(IF_ID__n561), .Y(IF_ID__n163) );
  BUFx6f_ASAP7_75t_R IF_ID___U303 ( .A(IF_ID__n165), .Y(IF_ID__n164) );
  BUFx6f_ASAP7_75t_R IF_ID___U304 ( .A(IF_ID__n167), .Y(IF_ID__n166) );
  BUFx6f_ASAP7_75t_R IF_ID___U305 ( .A(IF_ID__n169), .Y(IF_ID__n168) );
  BUFx2_ASAP7_75t_R IF_ID___U306 ( .A(IF_ID__n593), .Y(IF_ID__n172) );
  INVx3_ASAP7_75t_R IF_ID___U307 ( .A(IF_ID__n186), .Y(IF_ID__n357) );
  BUFx2_ASAP7_75t_R IF_ID___U308 ( .A(IF_ID__n665), .Y(IF_ID__n174) );
  BUFx2_ASAP7_75t_R IF_ID___U309 ( .A(IF_ID__n176), .Y(IF_ID__n175) );
  INVx1_ASAP7_75t_R IF_ID___U310 ( .A(IF_ID__n101), .Y(IF_ID__n177) );
  INVx1_ASAP7_75t_R IF_ID___U311 ( .A(IF_ID__n107), .Y(IF_ID__n179) );
  INVx1_ASAP7_75t_R IF_ID___U312 ( .A(IF_ID__n81), .Y(IF_ID__n181) );
  AO22x1_ASAP7_75t_R IF_ID___U313 ( .A1(inst_addr_o[15]), .A2(IF_ID__n31), .B1(
        IF_ID_inst_addr[15]), .B2(IF_ID__n513), .Y(IF_ID__n609) );
  INVx1_ASAP7_75t_R IF_ID___U314 ( .A(IF_ID__n97), .Y(IF_ID__n183) );
  BUFx4f_ASAP7_75t_R IF_ID___U315 ( .A(IF_ID__n479), .Y(IF_ID_inst_addr[4]) );
  BUFx4f_ASAP7_75t_R IF_ID___U316 ( .A(IF_ID__n588), .Y(IF_ID__n184) );
  BUFx4f_ASAP7_75t_R IF_ID___U317 ( .A(IF_ID__n563), .Y(IF_ID__n185) );
  BUFx6f_ASAP7_75t_R IF_ID___U318 ( .A(IF_ID__n187), .Y(IF_ID__n186) );
  BUFx6f_ASAP7_75t_R IF_ID___U319 ( .A(IF_ID__n189), .Y(IF_ID__n188) );
  BUFx4f_ASAP7_75t_R IF_ID___U320 ( .A(IF_ID__n566), .Y(IF_ID__n189) );
  INVx1_ASAP7_75t_R IF_ID___U321 ( .A(IF_ID__n157), .Y(IF_ID__n190) );
  BUFx2_ASAP7_75t_R IF_ID___U322 ( .A(IF_ID__n631), .Y(IF_ID__n191) );
  BUFx2_ASAP7_75t_R IF_ID___U323 ( .A(IF_ID__n634), .Y(IF_ID__n192) );
  BUFx2_ASAP7_75t_R IF_ID___U324 ( .A(IF_ID__n552), .Y(IF_ID__n193) );
  BUFx2_ASAP7_75t_R IF_ID___U325 ( .A(IF_ID__n550), .Y(IF_ID__n194) );
  BUFx2_ASAP7_75t_R IF_ID___U326 ( .A(IF_ID__n549), .Y(IF_ID__n195) );
  BUFx2_ASAP7_75t_R IF_ID___U327 ( .A(IF_ID__n639), .Y(IF_ID__n196) );
  BUFx5_ASAP7_75t_R IF_ID___U328 ( .A(IF_ID__n674), .Y(IF_ID__n249) );
  BUFx2_ASAP7_75t_R IF_ID___U329 ( .A(IF_ID__n661), .Y(IF_ID__n197) );
  BUFx2_ASAP7_75t_R IF_ID___U330 ( .A(IF_ID__n581), .Y(IF_ID__n198) );
  BUFx2_ASAP7_75t_R IF_ID___U331 ( .A(IF_ID__n666), .Y(IF_ID__n199) );
  BUFx2_ASAP7_75t_R IF_ID___U332 ( .A(IF_ID__n571), .Y(IF_ID__n200) );
  BUFx12f_ASAP7_75t_R IF_ID___U333 ( .A(IF_ID__n413), .Y(IF_ID_inst[24]) );
  BUFx3_ASAP7_75t_R IF_ID___U334 ( .A(IF_ID__n202), .Y(IF_ID__n201) );
  BUFx2_ASAP7_75t_R IF_ID___U335 ( .A(IF_ID__n676), .Y(IF_ID__n202) );
  AO22x1_ASAP7_75t_R IF_ID___U336 ( .A1(inst_addr_o[14]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[14]), .B2(IF_ID__n513), .Y(IF_ID__n610) );
  INVx1_ASAP7_75t_R IF_ID___U337 ( .A(IF_ID__n109), .Y(IF_ID__n205) );
  AO22x1_ASAP7_75t_R IF_ID___U338 ( .A1(inst_addr_o[8]), .A2(IF_ID__n21), .B1(
        IF_ID_inst_addr[8]), .B2(IF_ID__n516), .Y(IF_ID__n616) );
  INVx1_ASAP7_75t_R IF_ID___U339 ( .A(IF_ID__n105), .Y(IF_ID__n207) );
  AO22x1_ASAP7_75t_R IF_ID___U340 ( .A1(inst_addr_o[25]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[25]), .B2(IF_ID__n514), .Y(IF_ID__n601) );
  INVx6_ASAP7_75t_R IF_ID___U341 ( .A(IF_ID__n113), .Y(IF_ID__n514) );
  BUFx3_ASAP7_75t_R IF_ID___U342 ( .A(IF_ID__n211), .Y(IF_ID__n210) );
  BUFx2_ASAP7_75t_R IF_ID___U343 ( .A(IF_ID__n677), .Y(IF_ID__n211) );
  BUFx12f_ASAP7_75t_R IF_ID___U344 ( .A(IF_ID__n533), .Y(IF_ID__n215) );
  BUFx12f_ASAP7_75t_R IF_ID___U345 ( .A(IF_ID__n515), .Y(IF_ID__n533) );
  BUFx4f_ASAP7_75t_R IF_ID___U346 ( .A(IF_ID__n455), .Y(IF_ID_inst_addr[17]) );
  BUFx4f_ASAP7_75t_R IF_ID___U347 ( .A(IF_ID__n435), .Y(IF_ID_inst_addr[12]) );
  BUFx6f_ASAP7_75t_R IF_ID___U348 ( .A(IF_ID__n218), .Y(IF_ID__n217) );
  BUFx6f_ASAP7_75t_R IF_ID___U349 ( .A(IF_ID__n220), .Y(IF_ID__n219) );
  BUFx4f_ASAP7_75t_R IF_ID___U350 ( .A(IF_ID__n569), .Y(IF_ID__n220) );
  BUFx6f_ASAP7_75t_R IF_ID___U351 ( .A(IF_ID__n224), .Y(IF_ID__n223) );
  BUFx4f_ASAP7_75t_R IF_ID___U352 ( .A(IF_ID__n587), .Y(IF_ID__n224) );
  BUFx6f_ASAP7_75t_R IF_ID___U353 ( .A(IF_ID__n385), .Y(IF_ID_inst_addr[20]) );
  BUFx6f_ASAP7_75t_R IF_ID___U354 ( .A(IF_ID__n481), .Y(IF_ID_inst_addr[3]) );
  BUFx12f_ASAP7_75t_R IF_ID___U355 ( .A(IF_ID__n226), .Y(IF_ID__n225) );
  BUFx12f_ASAP7_75t_R IF_ID___U356 ( .A(IF_ID__n425), .Y(IF_ID__n226) );
  BUFx12f_ASAP7_75t_R IF_ID___U357 ( .A(IF_ID__n326), .Y(IF_ID__n227) );
  INVx2_ASAP7_75t_R IF_ID___U358 ( .A(IF_ID_opcode[6]), .Y(IF_ID__n235) );
  BUFx3_ASAP7_75t_R IF_ID___U359 ( .A(IF_ID__n747), .Y(IF_ID__n228) );
  INVx1_ASAP7_75t_R IF_ID___U360 ( .A(IF_ID__n146), .Y(IF_ID__n229) );
  INVx1_ASAP7_75t_R IF_ID___U361 ( .A(IF_ID__n148), .Y(IF_ID__n230) );
  INVx1_ASAP7_75t_R IF_ID___U362 ( .A(IF_ID__n86), .Y(IF_ID__n231) );
  AO22x1_ASAP7_75t_R IF_ID___U363 ( .A1(inst_addr_o[13]), .A2(IF_ID__n4), .B1(
        IF_ID_inst_addr[13]), .B2(IF_ID__n518), .Y(IF_ID__n611) );
  BUFx2_ASAP7_75t_R IF_ID___U364 ( .A(IF_ID__n594), .Y(IF_ID__n232) );
  BUFx2_ASAP7_75t_R IF_ID___U365 ( .A(IF_ID__n633), .Y(IF_ID__n233) );
  BUFx2_ASAP7_75t_R IF_ID___U366 ( .A(IF_ID__n635), .Y(IF_ID__n234) );
  BUFx5_ASAP7_75t_R IF_ID___U367 ( .A(IF_ID__n672), .Y(IF_ID__n326) );
  INVx2_ASAP7_75t_R IF_ID___U368 ( .A(IF_ID_opcode[5]), .Y(IF_ID__n589) );
  BUFx2_ASAP7_75t_R IF_ID___U369 ( .A(IF_ID__n660), .Y(IF_ID__n236) );
  BUFx2_ASAP7_75t_R IF_ID___U370 ( .A(IF_ID__n583), .Y(IF_ID__n237) );
  BUFx2_ASAP7_75t_R IF_ID___U371 ( .A(IF_ID__n662), .Y(IF_ID__n238) );
  INVx2_ASAP7_75t_R IF_ID___U372 ( .A(IF_ID__n518), .Y(IF_ID__n530) );
  BUFx12f_ASAP7_75t_R IF_ID___U373 ( .A(IF_ID__n421), .Y(IF_ID_inst[14]) );
  BUFx6f_ASAP7_75t_R IF_ID___U374 ( .A(IF_ID__n457), .Y(IF_ID_inst_addr[16]) );
  BUFx3_ASAP7_75t_R IF_ID___U375 ( .A(IF_ID__n243), .Y(IF_ID__n242) );
  BUFx2_ASAP7_75t_R IF_ID___U376 ( .A(IF_ID__n729), .Y(IF_ID__n243) );
  BUFx2_ASAP7_75t_R IF_ID___U377 ( .A(IF_ID__n591), .Y(IF_ID__n244) );
  BUFx2_ASAP7_75t_R IF_ID___U378 ( .A(IF_ID__n670), .Y(IF_ID__n247) );
  BUFx6f_ASAP7_75t_R IF_ID___U379 ( .A(IF_ID__n251), .Y(IF_ID__n250) );
  BUFx4f_ASAP7_75t_R IF_ID___U380 ( .A(IF_ID__n228), .Y(IF_ID__n251) );
  BUFx12f_ASAP7_75t_R IF_ID___U381 ( .A(IF_ID__n329), .Y(IF_ID_inst[27]) );
  BUFx6f_ASAP7_75t_R IF_ID___U382 ( .A(IF_ID__n387), .Y(IF_ID_inst_addr[1]) );
  BUFx2_ASAP7_75t_R IF_ID___U383 ( .A(IF_ID__n254), .Y(IF_ID__n252) );
  BUFx6f_ASAP7_75t_R IF_ID___U384 ( .A(IF_ID__n254), .Y(IF_ID_inst_addr[6]) );
  BUFx6f_ASAP7_75t_R IF_ID___U385 ( .A(IF_ID__n474), .Y(IF_ID__n254) );
  BUFx4f_ASAP7_75t_R IF_ID___U386 ( .A(IF_ID__n475), .Y(IF_ID__n474) );
  BUFx3_ASAP7_75t_R IF_ID___U387 ( .A(IF_ID__n339), .Y(IF_ID__n475) );
  BUFx4f_ASAP7_75t_R IF_ID___U388 ( .A(IF_ID__n308), .Y(IF_ID__n389) );
  BUFx3_ASAP7_75t_R IF_ID___U389 ( .A(IF_ID__n256), .Y(IF_ID__n255) );
  BUFx2_ASAP7_75t_R IF_ID___U390 ( .A(IF_ID__n725), .Y(IF_ID__n256) );
  BUFx3_ASAP7_75t_R IF_ID___U391 ( .A(IF_ID__n258), .Y(IF_ID__n257) );
  BUFx2_ASAP7_75t_R IF_ID___U392 ( .A(IF_ID__n726), .Y(IF_ID__n258) );
  BUFx3_ASAP7_75t_R IF_ID___U393 ( .A(IF_ID__n260), .Y(IF_ID__n259) );
  BUFx2_ASAP7_75t_R IF_ID___U394 ( .A(IF_ID__n728), .Y(IF_ID__n260) );
  BUFx12f_ASAP7_75t_R IF_ID___U395 ( .A(IF_ID__n262), .Y(IF_ID__n261) );
  BUFx12f_ASAP7_75t_R IF_ID___U396 ( .A(IF_ID__n417), .Y(IF_ID__n262) );
  BUFx3_ASAP7_75t_R IF_ID___U397 ( .A(IF_ID__n264), .Y(IF_ID__n263) );
  BUFx2_ASAP7_75t_R IF_ID___U398 ( .A(IF_ID__n736), .Y(IF_ID__n264) );
  BUFx3_ASAP7_75t_R IF_ID___U399 ( .A(IF_ID__n266), .Y(IF_ID__n265) );
  BUFx2_ASAP7_75t_R IF_ID___U400 ( .A(IF_ID__n742), .Y(IF_ID__n266) );
  BUFx12f_ASAP7_75t_R IF_ID___U401 ( .A(IF_ID__n268), .Y(IF_ID__n267) );
  BUFx12f_ASAP7_75t_R IF_ID___U402 ( .A(IF_ID__n500), .Y(IF_ID__n268) );
  BUFx2_ASAP7_75t_R IF_ID___U403 ( .A(IF_ID__n592), .Y(IF_ID__n269) );
  BUFx2_ASAP7_75t_R IF_ID___U404 ( .A(IF_ID__n557), .Y(IF_ID__n270) );
  BUFx6f_ASAP7_75t_R IF_ID___U405 ( .A(IF_ID__n437), .Y(IF_ID_inst_addr[31]) );
  BUFx6f_ASAP7_75t_R IF_ID___U406 ( .A(IF_ID__n441), .Y(IF_ID_inst_addr[26]) );
  BUFx6f_ASAP7_75t_R IF_ID___U407 ( .A(IF_ID__n389), .Y(IF_ID_inst_addr[0]) );
  BUFx6f_ASAP7_75t_R IF_ID___U408 ( .A(IF_ID__n483), .Y(IF_ID_rd[4]) );
  BUFx6f_ASAP7_75t_R IF_ID___U409 ( .A(IF_ID__n489), .Y(IF_ID_rd[1]) );
  BUFx4f_ASAP7_75t_R IF_ID___U410 ( .A(IF_ID__n340), .Y(IF_ID__n391) );
  BUFx4f_ASAP7_75t_R IF_ID___U411 ( .A(IF_ID__n380), .Y(IF_ID__n443) );
  BUFx4f_ASAP7_75t_R IF_ID___U412 ( .A(IF_ID__n381), .Y(IF_ID__n451) );
  BUFx4f_ASAP7_75t_R IF_ID___U413 ( .A(IF_ID__n343), .Y(IF_ID__n399) );
  BUFx4f_ASAP7_75t_R IF_ID___U414 ( .A(IF_ID__n485), .Y(IF_ID_rd[3]) );
  BUFx4f_ASAP7_75t_R IF_ID___U415 ( .A(IF_ID__n491), .Y(IF_ID_rd[0]) );
  BUFx3_ASAP7_75t_R IF_ID___U416 ( .A(IF_ID__n272), .Y(IF_ID__n271) );
  BUFx2_ASAP7_75t_R IF_ID___U417 ( .A(IF_ID__n721), .Y(IF_ID__n272) );
  BUFx3_ASAP7_75t_R IF_ID___U418 ( .A(IF_ID__n274), .Y(IF_ID__n273) );
  BUFx2_ASAP7_75t_R IF_ID___U419 ( .A(IF_ID__n723), .Y(IF_ID__n274) );
  BUFx3_ASAP7_75t_R IF_ID___U420 ( .A(IF_ID__n276), .Y(IF_ID__n275) );
  BUFx2_ASAP7_75t_R IF_ID___U421 ( .A(IF_ID__n724), .Y(IF_ID__n276) );
  BUFx3_ASAP7_75t_R IF_ID___U422 ( .A(IF_ID__n278), .Y(IF_ID__n277) );
  BUFx2_ASAP7_75t_R IF_ID___U423 ( .A(IF_ID__n727), .Y(IF_ID__n278) );
  BUFx12f_ASAP7_75t_R IF_ID___U424 ( .A(IF_ID__n280), .Y(IF_ID__n279) );
  BUFx12f_ASAP7_75t_R IF_ID___U425 ( .A(IF_ID__n415), .Y(IF_ID__n280) );
  BUFx3_ASAP7_75t_R IF_ID___U426 ( .A(IF_ID__n282), .Y(IF_ID__n281) );
  BUFx2_ASAP7_75t_R IF_ID___U427 ( .A(IF_ID__n731), .Y(IF_ID__n282) );
  BUFx3_ASAP7_75t_R IF_ID___U428 ( .A(IF_ID__n284), .Y(IF_ID__n283) );
  BUFx2_ASAP7_75t_R IF_ID___U429 ( .A(IF_ID__n732), .Y(IF_ID__n284) );
  BUFx3_ASAP7_75t_R IF_ID___U430 ( .A(IF_ID__n286), .Y(IF_ID__n285) );
  BUFx2_ASAP7_75t_R IF_ID___U431 ( .A(IF_ID__n733), .Y(IF_ID__n286) );
  BUFx3_ASAP7_75t_R IF_ID___U432 ( .A(IF_ID__n288), .Y(IF_ID__n287) );
  BUFx2_ASAP7_75t_R IF_ID___U433 ( .A(IF_ID__n734), .Y(IF_ID__n288) );
  BUFx3_ASAP7_75t_R IF_ID___U434 ( .A(IF_ID__n290), .Y(IF_ID__n289) );
  BUFx2_ASAP7_75t_R IF_ID___U435 ( .A(IF_ID__n735), .Y(IF_ID__n290) );
  BUFx3_ASAP7_75t_R IF_ID___U436 ( .A(IF_ID__n292), .Y(IF_ID__n291) );
  BUFx2_ASAP7_75t_R IF_ID___U437 ( .A(IF_ID__n739), .Y(IF_ID__n292) );
  BUFx3_ASAP7_75t_R IF_ID___U438 ( .A(IF_ID__n294), .Y(IF_ID__n293) );
  BUFx2_ASAP7_75t_R IF_ID___U439 ( .A(IF_ID__n741), .Y(IF_ID__n294) );
  OR2x2_ASAP7_75t_R IF_ID___U440 ( .A(IF_ID__n295), .B(IF_ID__n520), .Y(IF_ID__n671) );
  OR2x2_ASAP7_75t_R IF_ID___U441 ( .A(IF_ID__n529), .B(IF_ID__n564), .Y(IF_ID__n519) );
  INVx1_ASAP7_75t_R IF_ID___U442 ( .A(IF_ID__n162), .Y(IF_ID__n295) );
  BUFx6f_ASAP7_75t_R IF_ID___U443 ( .A(IF_ID__n391), .Y(IF_ID_inst_addr[30]) );
  BUFx6f_ASAP7_75t_R IF_ID___U444 ( .A(IF_ID__n443), .Y(IF_ID_inst_addr[24]) );
  BUFx6f_ASAP7_75t_R IF_ID___U445 ( .A(IF_ID__n451), .Y(IF_ID_inst_addr[19]) );
  BUFx6f_ASAP7_75t_R IF_ID___U446 ( .A(IF_ID__n399), .Y(IF_ID_inst_addr[2]) );
  BUFx12f_ASAP7_75t_R IF_ID___U447 ( .A(IF_ID__n279), .Y(IF_ID_inst[23]) );
  BUFx12f_ASAP7_75t_R IF_ID___U448 ( .A(IF_ID__n225), .Y(IF_ID_inst[17]) );
  BUFx12f_ASAP7_75t_R IF_ID___U449 ( .A(IF_ID__n494), .Y(IF_ID_inst[11]) );
  BUFx2_ASAP7_75t_R IF_ID___U450 ( .A(IF_ID__n697), .Y(IF_ID__n300) );
  BUFx2_ASAP7_75t_R IF_ID___U451 ( .A(IF_ID__n701), .Y(IF_ID__n301) );
  BUFx2_ASAP7_75t_R IF_ID___U452 ( .A(IF_ID__n704), .Y(IF_ID__n302) );
  BUFx2_ASAP7_75t_R IF_ID___U453 ( .A(IF_ID__n706), .Y(IF_ID__n303) );
  BUFx2_ASAP7_75t_R IF_ID___U454 ( .A(IF_ID__n708), .Y(IF_ID__n304) );
  BUFx2_ASAP7_75t_R IF_ID___U455 ( .A(IF_ID__n715), .Y(IF_ID__n306) );
  BUFx2_ASAP7_75t_R IF_ID___U456 ( .A(IF_ID__n717), .Y(IF_ID__n307) );
  BUFx2_ASAP7_75t_R IF_ID___U457 ( .A(IF_ID__n718), .Y(IF_ID__n308) );
  BUFx3_ASAP7_75t_R IF_ID___U458 ( .A(IF_ID__n310), .Y(IF_ID__n309) );
  BUFx2_ASAP7_75t_R IF_ID___U459 ( .A(IF_ID__n680), .Y(IF_ID__n310) );
  BUFx4f_ASAP7_75t_R IF_ID___U460 ( .A(IF_ID__n309), .Y(IF_ID__n487) );
  BUFx3_ASAP7_75t_R IF_ID___U461 ( .A(IF_ID__n312), .Y(IF_ID__n311) );
  BUFx2_ASAP7_75t_R IF_ID___U462 ( .A(IF_ID__n720), .Y(IF_ID__n312) );
  BUFx3_ASAP7_75t_R IF_ID___U463 ( .A(IF_ID__n314), .Y(IF_ID__n313) );
  BUFx2_ASAP7_75t_R IF_ID___U464 ( .A(IF_ID__n722), .Y(IF_ID__n314) );
  BUFx3_ASAP7_75t_R IF_ID___U465 ( .A(IF_ID__n316), .Y(IF_ID__n315) );
  BUFx2_ASAP7_75t_R IF_ID___U466 ( .A(IF_ID__n738), .Y(IF_ID__n316) );
  BUFx3_ASAP7_75t_R IF_ID___U467 ( .A(IF_ID__n318), .Y(IF_ID__n317) );
  BUFx2_ASAP7_75t_R IF_ID___U468 ( .A(IF_ID__n740), .Y(IF_ID__n318) );
  INVx1_ASAP7_75t_R IF_ID___U469 ( .A(IF_ID__n129), .Y(IF_ID__n320) );
  INVx1_ASAP7_75t_R IF_ID___U470 ( .A(IF_ID__n96), .Y(IF_ID__n321) );
  AO22x1_ASAP7_75t_R IF_ID___U471 ( .A1(inst_addr_o[9]), .A2(IF_ID__n21), .B1(
        IF_ID_inst_addr[9]), .B2(IF_ID__n515), .Y(IF_ID__n615) );
  INVx1_ASAP7_75t_R IF_ID___U472 ( .A(IF_ID__n133), .Y(IF_ID__n322) );
  AO22x1_ASAP7_75t_R IF_ID___U473 ( .A1(inst_addr_o[28]), .A2(IF_ID__n28), .B1(
        IF_ID_inst_addr[28]), .B2(IF_ID__n515), .Y(IF_ID__n598) );
  INVx1_ASAP7_75t_R IF_ID___U474 ( .A(IF_ID__n175), .Y(IF_ID__n323) );
  BUFx4f_ASAP7_75t_R IF_ID___U475 ( .A(IF_ID__n325), .Y(IF_ID__n324) );
  INVx2_ASAP7_75t_R IF_ID___U476 ( .A(IF_ID__n185), .Y(IF_ID__n325) );
  INVx1_ASAP7_75t_R IF_ID___U477 ( .A(IF_ID__n324), .Y(IF_ID__n520) );
  BUFx4f_ASAP7_75t_R IF_ID___U478 ( .A(IF_ID__n273), .Y(IF_ID__n329) );
  BUFx6f_ASAP7_75t_R IF_ID___U479 ( .A(IF_ID__n331), .Y(IF_ID_inst[26]) );
  BUFx4f_ASAP7_75t_R IF_ID___U480 ( .A(IF_ID__n275), .Y(IF_ID__n331) );
  BUFx6f_ASAP7_75t_R IF_ID___U481 ( .A(IF_ID__n333), .Y(IF_ID_inst[25]) );
  BUFx4f_ASAP7_75t_R IF_ID___U482 ( .A(IF_ID__n255), .Y(IF_ID__n333) );
  BUFx6f_ASAP7_75t_R IF_ID___U483 ( .A(IF_ID__n335), .Y(IF_ID_opcode[1]) );
  BUFx4f_ASAP7_75t_R IF_ID___U484 ( .A(IF_ID__n201), .Y(IF_ID__n335) );
  BUFx2_ASAP7_75t_R IF_ID___U485 ( .A(IF_ID__n640), .Y(IF_ID__n336) );
  BUFx2_ASAP7_75t_R IF_ID___U486 ( .A(IF_ID__n546), .Y(IF_ID__n337) );
  BUFx6f_ASAP7_75t_R IF_ID___U487 ( .A(IF_ID__n487), .Y(IF_ID_rd[2]) );
  BUFx12f_ASAP7_75t_R IF_ID___U488 ( .A(IF_ID__n261), .Y(IF_ID_inst[22]) );
  BUFx12f_ASAP7_75t_R IF_ID___U489 ( .A(IF_ID__n427), .Y(IF_ID_inst[16]) );
  BUFx12f_ASAP7_75t_R IF_ID___U490 ( .A(IF_ID__n496), .Y(IF_ID_inst[10]) );
  BUFx12f_ASAP7_75t_R IF_ID___U491 ( .A(IF_ID__n267), .Y(IF_ID_inst[8]) );
  BUFx2_ASAP7_75t_R IF_ID___U492 ( .A(IF_ID__n710), .Y(IF_ID__n338) );
  BUFx2_ASAP7_75t_R IF_ID___U493 ( .A(IF_ID__n712), .Y(IF_ID__n339) );
  BUFx2_ASAP7_75t_R IF_ID___U494 ( .A(IF_ID__n688), .Y(IF_ID__n340) );
  BUFx2_ASAP7_75t_R IF_ID___U495 ( .A(IF_ID__n698), .Y(IF_ID__n341) );
  BUFx2_ASAP7_75t_R IF_ID___U496 ( .A(IF_ID__n702), .Y(IF_ID__n342) );
  BUFx2_ASAP7_75t_R IF_ID___U497 ( .A(IF_ID__n716), .Y(IF_ID__n343) );
  BUFx2_ASAP7_75t_R IF_ID___U498 ( .A(IF_ID__n678), .Y(IF_ID__n344) );
  BUFx2_ASAP7_75t_R IF_ID___U499 ( .A(IF_ID__n679), .Y(IF_ID__n345) );
  BUFx2_ASAP7_75t_R IF_ID___U500 ( .A(IF_ID__n681), .Y(IF_ID__n346) );
  BUFx2_ASAP7_75t_R IF_ID___U501 ( .A(IF_ID__n682), .Y(IF_ID__n347) );
  BUFx3_ASAP7_75t_R IF_ID___U502 ( .A(IF_ID__n349), .Y(IF_ID__n348) );
  BUFx2_ASAP7_75t_R IF_ID___U503 ( .A(IF_ID__n737), .Y(IF_ID__n349) );
  BUFx3_ASAP7_75t_R IF_ID___U504 ( .A(IF_ID__n351), .Y(IF_ID__n350) );
  BUFx2_ASAP7_75t_R IF_ID___U505 ( .A(IF_ID__n743), .Y(IF_ID__n351) );
  BUFx12f_ASAP7_75t_R IF_ID___U506 ( .A(IF_ID__n353), .Y(IF_ID__n352) );
  BUFx12f_ASAP7_75t_R IF_ID___U507 ( .A(IF_ID__n502), .Y(IF_ID__n353) );
  AO22x1_ASAP7_75t_R IF_ID___U508 ( .A1(inst_addr_o[29]), .A2(IF_ID__n21), .B1(
        IF_ID_inst_addr[29]), .B2(IF_ID__n518), .Y(IF_ID__n597) );
  BUFx12f_ASAP7_75t_R IF_ID___U509 ( .A(IF_ID__n730), .Y(IF_ID__n355) );
  AND2x4_ASAP7_75t_R IF_ID___U510 ( .A(inst_i[16]), .B(IF_ID__n30), .Y(IF_ID__n565) );
  BUFx6f_ASAP7_75t_R IF_ID___U511 ( .A(IF_ID__n365), .Y(IF_ID_inst[30]) );
  BUFx4f_ASAP7_75t_R IF_ID___U512 ( .A(IF_ID__n311), .Y(IF_ID__n365) );
  BUFx6f_ASAP7_75t_R IF_ID___U513 ( .A(IF_ID__n367), .Y(IF_ID_inst[29]) );
  BUFx4f_ASAP7_75t_R IF_ID___U514 ( .A(IF_ID__n271), .Y(IF_ID__n367) );
  BUFx6f_ASAP7_75t_R IF_ID___U515 ( .A(IF_ID__n369), .Y(IF_ID_inst[28]) );
  BUFx4f_ASAP7_75t_R IF_ID___U516 ( .A(IF_ID__n313), .Y(IF_ID__n369) );
  BUFx6f_ASAP7_75t_R IF_ID___U517 ( .A(IF_ID__n371), .Y(IF_ID_inst[19]) );
  BUFx4f_ASAP7_75t_R IF_ID___U518 ( .A(IF_ID__n281), .Y(IF_ID__n371) );
  BUFx6f_ASAP7_75t_R IF_ID___U519 ( .A(IF_ID__n373), .Y(IF_ID_inst[18]) );
  BUFx4f_ASAP7_75t_R IF_ID___U520 ( .A(IF_ID__n283), .Y(IF_ID__n373) );
  BUFx12f_ASAP7_75t_R IF_ID___U521 ( .A(IF_ID__n375), .Y(IF_ID_inst[5]) );
  BUFx12f_ASAP7_75t_R IF_ID___U522 ( .A(IF_ID__n498), .Y(IF_ID_inst[9]) );
  BUFx12f_ASAP7_75t_R IF_ID___U523 ( .A(IF_ID__n352), .Y(IF_ID_inst[7]) );
  BUFx4f_ASAP7_75t_R IF_ID___U524 ( .A(IF_ID__n377), .Y(IF_ID__n376) );
  INVx2_ASAP7_75t_R IF_ID___U525 ( .A(IF_ID__n184), .Y(IF_ID__n377) );
  BUFx2_ASAP7_75t_R IF_ID___U526 ( .A(IF_ID__n687), .Y(IF_ID__n378) );
  BUFx2_ASAP7_75t_R IF_ID___U527 ( .A(IF_ID__n692), .Y(IF_ID__n379) );
  BUFx2_ASAP7_75t_R IF_ID___U528 ( .A(IF_ID__n694), .Y(IF_ID__n380) );
  BUFx2_ASAP7_75t_R IF_ID___U529 ( .A(IF_ID__n699), .Y(IF_ID__n381) );
  INVx1_ASAP7_75t_R IF_ID___U530 ( .A(IF_ID__n88), .Y(IF_ID__n382) );
  AO22x1_ASAP7_75t_R IF_ID___U531 ( .A1(inst_i[30]), .A2(IF_ID__n29), .B1(IF_ID_inst[30]), 
        .B2(IF_ID__n13), .Y(IF_ID__n625) );
  INVx1_ASAP7_75t_R IF_ID___U532 ( .A(IF_ID__n152), .Y(IF_ID__n383) );
  BUFx3_ASAP7_75t_R IF_ID___U533 ( .A(IF_ID__n341), .Y(IF_ID__n385) );
  BUFx3_ASAP7_75t_R IF_ID___U534 ( .A(IF_ID__n307), .Y(IF_ID__n387) );
  BUFx3_ASAP7_75t_R IF_ID___U535 ( .A(IF_ID__n393), .Y(IF_ID_inst_addr[29]) );
  BUFx2_ASAP7_75t_R IF_ID___U536 ( .A(IF_ID__n689), .Y(IF_ID__n393) );
  BUFx3_ASAP7_75t_R IF_ID___U537 ( .A(IF_ID__n395), .Y(IF_ID_inst_addr[28]) );
  BUFx2_ASAP7_75t_R IF_ID___U538 ( .A(IF_ID__n690), .Y(IF_ID__n395) );
  BUFx3_ASAP7_75t_R IF_ID___U539 ( .A(IF_ID__n397), .Y(IF_ID_inst_addr[25]) );
  BUFx2_ASAP7_75t_R IF_ID___U540 ( .A(IF_ID__n693), .Y(IF_ID__n397) );
  INVx2_ASAP7_75t_R IF_ID___U541 ( .A(IF_ID__n578), .Y(IF_ID__n401) );
  BUFx6f_ASAP7_75t_R IF_ID___U542 ( .A(IF_ID__n409), .Y(IF_ID_inst[13]) );
  BUFx4f_ASAP7_75t_R IF_ID___U543 ( .A(IF_ID__n348), .Y(IF_ID__n409) );
  BUFx6f_ASAP7_75t_R IF_ID___U544 ( .A(IF_ID__n411), .Y(IF_ID_opcode[0]) );
  BUFx4f_ASAP7_75t_R IF_ID___U545 ( .A(IF_ID__n210), .Y(IF_ID__n411) );
  BUFx4f_ASAP7_75t_R IF_ID___U546 ( .A(IF_ID__n257), .Y(IF_ID__n413) );
  BUFx4f_ASAP7_75t_R IF_ID___U547 ( .A(IF_ID__n277), .Y(IF_ID__n415) );
  BUFx4f_ASAP7_75t_R IF_ID___U548 ( .A(IF_ID__n259), .Y(IF_ID__n417) );
  BUFx6f_ASAP7_75t_R IF_ID___U549 ( .A(IF_ID__n419), .Y(IF_ID_inst[21]) );
  BUFx4f_ASAP7_75t_R IF_ID___U550 ( .A(IF_ID__n242), .Y(IF_ID__n419) );
  BUFx4f_ASAP7_75t_R IF_ID___U551 ( .A(IF_ID__n263), .Y(IF_ID__n421) );
  BUFx6f_ASAP7_75t_R IF_ID___U552 ( .A(IF_ID__n423), .Y(IF_ID_inst[12]) );
  BUFx4f_ASAP7_75t_R IF_ID___U553 ( .A(IF_ID__n315), .Y(IF_ID__n423) );
  BUFx4f_ASAP7_75t_R IF_ID___U554 ( .A(IF_ID__n285), .Y(IF_ID__n425) );
  BUFx4f_ASAP7_75t_R IF_ID___U555 ( .A(IF_ID__n287), .Y(IF_ID__n427) );
  BUFx6f_ASAP7_75t_R IF_ID___U556 ( .A(IF_ID__n429), .Y(IF_ID_inst[15]) );
  BUFx4f_ASAP7_75t_R IF_ID___U557 ( .A(IF_ID__n289), .Y(IF_ID__n429) );
  BUFx12f_ASAP7_75t_R IF_ID___U558 ( .A(IF_ID__n431), .Y(IF_ID_opcode[6]) );
  BUFx12f_ASAP7_75t_R IF_ID___U559 ( .A(IF_ID__n227), .Y(IF_ID__n431) );
  BUFx2_ASAP7_75t_R IF_ID___U560 ( .A(IF_ID__n303), .Y(IF_ID__n435) );
  BUFx3_ASAP7_75t_R IF_ID___U561 ( .A(IF_ID__n378), .Y(IF_ID__n437) );
  BUFx3_ASAP7_75t_R IF_ID___U562 ( .A(IF_ID__n439), .Y(IF_ID_inst_addr[27]) );
  BUFx2_ASAP7_75t_R IF_ID___U563 ( .A(IF_ID__n691), .Y(IF_ID__n439) );
  BUFx3_ASAP7_75t_R IF_ID___U564 ( .A(IF_ID__n379), .Y(IF_ID__n441) );
  BUFx3_ASAP7_75t_R IF_ID___U565 ( .A(IF_ID__n445), .Y(IF_ID_inst_addr[23]) );
  BUFx2_ASAP7_75t_R IF_ID___U566 ( .A(IF_ID__n695), .Y(IF_ID__n445) );
  BUFx2_ASAP7_75t_R IF_ID___U567 ( .A(IF_ID__n696), .Y(IF_ID__n447) );
  BUFx3_ASAP7_75t_R IF_ID___U568 ( .A(IF_ID__n449), .Y(IF_ID_inst_addr[21]) );
  BUFx2_ASAP7_75t_R IF_ID___U569 ( .A(IF_ID__n300), .Y(IF_ID__n449) );
  BUFx2_ASAP7_75t_R IF_ID___U570 ( .A(IF_ID__n700), .Y(IF_ID__n453) );
  BUFx2_ASAP7_75t_R IF_ID___U571 ( .A(IF_ID__n301), .Y(IF_ID__n455) );
  BUFx3_ASAP7_75t_R IF_ID___U572 ( .A(IF_ID__n342), .Y(IF_ID__n457) );
  BUFx3_ASAP7_75t_R IF_ID___U573 ( .A(IF_ID__n459), .Y(IF_ID_inst_addr[15]) );
  BUFx2_ASAP7_75t_R IF_ID___U574 ( .A(IF_ID__n703), .Y(IF_ID__n459) );
  BUFx3_ASAP7_75t_R IF_ID___U575 ( .A(IF_ID__n461), .Y(IF_ID_inst_addr[14]) );
  BUFx2_ASAP7_75t_R IF_ID___U576 ( .A(IF_ID__n302), .Y(IF_ID__n461) );
  BUFx3_ASAP7_75t_R IF_ID___U577 ( .A(IF_ID__n463), .Y(IF_ID_inst_addr[13]) );
  BUFx2_ASAP7_75t_R IF_ID___U578 ( .A(IF_ID__n705), .Y(IF_ID__n463) );
  BUFx3_ASAP7_75t_R IF_ID___U579 ( .A(IF_ID__n465), .Y(IF_ID_inst_addr[11]) );
  BUFx2_ASAP7_75t_R IF_ID___U580 ( .A(IF_ID__n707), .Y(IF_ID__n465) );
  BUFx3_ASAP7_75t_R IF_ID___U581 ( .A(IF_ID__n467), .Y(IF_ID_inst_addr[10]) );
  BUFx2_ASAP7_75t_R IF_ID___U582 ( .A(IF_ID__n304), .Y(IF_ID__n467) );
  BUFx3_ASAP7_75t_R IF_ID___U583 ( .A(IF_ID__n469), .Y(IF_ID_inst_addr[9]) );
  BUFx2_ASAP7_75t_R IF_ID___U584 ( .A(IF_ID__n709), .Y(IF_ID__n469) );
  BUFx3_ASAP7_75t_R IF_ID___U585 ( .A(IF_ID__n471), .Y(IF_ID_inst_addr[8]) );
  BUFx2_ASAP7_75t_R IF_ID___U586 ( .A(IF_ID__n338), .Y(IF_ID__n471) );
  BUFx3_ASAP7_75t_R IF_ID___U587 ( .A(IF_ID__n473), .Y(IF_ID_inst_addr[7]) );
  BUFx2_ASAP7_75t_R IF_ID___U588 ( .A(IF_ID__n711), .Y(IF_ID__n473) );
  BUFx3_ASAP7_75t_R IF_ID___U589 ( .A(IF_ID__n477), .Y(IF_ID_inst_addr[5]) );
  BUFx2_ASAP7_75t_R IF_ID___U590 ( .A(IF_ID__n713), .Y(IF_ID__n477) );
  BUFx2_ASAP7_75t_R IF_ID___U591 ( .A(IF_ID__n714), .Y(IF_ID__n479) );
  BUFx3_ASAP7_75t_R IF_ID___U592 ( .A(IF_ID__n306), .Y(IF_ID__n481) );
  BUFx3_ASAP7_75t_R IF_ID___U593 ( .A(IF_ID__n344), .Y(IF_ID__n483) );
  BUFx3_ASAP7_75t_R IF_ID___U594 ( .A(IF_ID__n345), .Y(IF_ID__n485) );
  BUFx3_ASAP7_75t_R IF_ID___U595 ( .A(IF_ID__n346), .Y(IF_ID__n489) );
  BUFx3_ASAP7_75t_R IF_ID___U596 ( .A(IF_ID__n347), .Y(IF_ID__n491) );
  INVx2_ASAP7_75t_R IF_ID___U597 ( .A(IF_ID__n142), .Y(IF_ID__n492) );
  BUFx4f_ASAP7_75t_R IF_ID___U598 ( .A(IF_ID__n291), .Y(IF_ID__n494) );
  BUFx4f_ASAP7_75t_R IF_ID___U599 ( .A(IF_ID__n317), .Y(IF_ID__n496) );
  BUFx4f_ASAP7_75t_R IF_ID___U600 ( .A(IF_ID__n293), .Y(IF_ID__n498) );
  BUFx4f_ASAP7_75t_R IF_ID___U601 ( .A(IF_ID__n265), .Y(IF_ID__n500) );
  BUFx4f_ASAP7_75t_R IF_ID___U602 ( .A(IF_ID__n350), .Y(IF_ID__n502) );
  BUFx12f_ASAP7_75t_R IF_ID___U603 ( .A(IF_ID__n504), .Y(IF_ID_inst[20]) );
  BUFx12f_ASAP7_75t_R IF_ID___U604 ( .A(IF_ID__n355), .Y(IF_ID__n504) );
  BUFx12f_ASAP7_75t_R IF_ID___U605 ( .A(IF_ID__n506), .Y(IF_ID_opcode[4]) );
  BUFx12f_ASAP7_75t_R IF_ID___U606 ( .A(IF_ID__n249), .Y(IF_ID__n506) );
  BUFx12f_ASAP7_75t_R IF_ID___U607 ( .A(IF_ID__n508), .Y(IF_ID_opcode[5]) );
  BUFx12f_ASAP7_75t_R IF_ID___U608 ( .A(IF_ID__n673), .Y(IF_ID__n508) );
  BUFx12f_ASAP7_75t_R IF_ID___U609 ( .A(IF_ID__n510), .Y(IF_ID_inst[31]) );
  BUFx12f_ASAP7_75t_R IF_ID___U610 ( .A(IF_ID__n719), .Y(IF_ID__n510) );
  INVx1_ASAP7_75t_R IF_ID___U611 ( .A(IF_ID__n121), .Y(IF_ID__n535) );
  OA21x2_ASAP7_75t_R IF_ID___U612 ( .A1(IF_ID__n12), .A2(IF_ID__n118), .B(IF_ID__n141), .Y(IF_ID__n654) );
  INVx1_ASAP7_75t_R IF_ID___U613 ( .A(IF_ID__n139), .Y(IF_ID__n536) );
  OA21x2_ASAP7_75t_R IF_ID___U614 ( .A1(IF_ID__n12), .A2(IF_ID__n100), .B(IF_ID__n407), .Y(IF_ID__n653) );
  OA21x2_ASAP7_75t_R IF_ID___U615 ( .A1(IF_ID__n12), .A2(IF_ID__n537), .B(IF_ID__n406), .Y(IF_ID__n652) );
  OA21x2_ASAP7_75t_R IF_ID___U616 ( .A1(IF_ID__n12), .A2(IF_ID__n538), .B(IF_ID__n363), .Y(IF_ID__n651) );
  OA21x2_ASAP7_75t_R IF_ID___U617 ( .A1(IF_ID__n521), .A2(IF_ID__n539), .B(IF_ID__n405), .Y(IF_ID__n650) );
  OA21x2_ASAP7_75t_R IF_ID___U618 ( .A1(IF_ID__n521), .A2(IF_ID__n126), .B(IF_ID__n376), .Y(IF_ID__n649) );
  OA21x2_ASAP7_75t_R IF_ID___U619 ( .A1(IF_ID__n522), .A2(IF_ID__n190), .B(IF_ID__n362), .Y(IF_ID__n648) );
  OA21x2_ASAP7_75t_R IF_ID___U620 ( .A1(IF_ID__n541), .A2(IF_ID__n522), .B(IF_ID__n404), .Y(IF_ID__n647) );
  INVx1_ASAP7_75t_R IF_ID___U621 ( .A(IF_ID_inst[8]), .Y(IF_ID__n542) );
  OA21x2_ASAP7_75t_R IF_ID___U622 ( .A1(IF_ID__n523), .A2(IF_ID__n542), .B(IF_ID__n403), .Y(IF_ID__n646) );
  INVx1_ASAP7_75t_R IF_ID___U623 ( .A(IF_ID_inst[9]), .Y(IF_ID__n543) );
  OA21x2_ASAP7_75t_R IF_ID___U624 ( .A1(IF_ID__n523), .A2(IF_ID__n543), .B(IF_ID__n361), .Y(IF_ID__n645) );
  INVx1_ASAP7_75t_R IF_ID___U625 ( .A(IF_ID_inst[10]), .Y(IF_ID__n544) );
  OA21x2_ASAP7_75t_R IF_ID___U626 ( .A1(IF_ID__n524), .A2(IF_ID__n544), .B(IF_ID__n402), .Y(IF_ID__n644) );
  INVx1_ASAP7_75t_R IF_ID___U627 ( .A(IF_ID_inst[11]), .Y(IF_ID__n545) );
  OA21x2_ASAP7_75t_R IF_ID___U628 ( .A1(IF_ID__n524), .A2(IF_ID__n545), .B(IF_ID__n401), .Y(IF_ID__n643) );
  INVx1_ASAP7_75t_R IF_ID___U629 ( .A(IF_ID_inst[15]), .Y(IF_ID__n546) );
  OA21x2_ASAP7_75t_R IF_ID___U630 ( .A1(IF_ID__n527), .A2(IF_ID__n337), .B(IF_ID__n324), .Y(IF_ID__n640) );
  INVx1_ASAP7_75t_R IF_ID___U631 ( .A(IF_ID_inst[16]), .Y(IF_ID__n547) );
  OA21x2_ASAP7_75t_R IF_ID___U632 ( .A1(IF_ID__n527), .A2(IF_ID__n547), .B(IF_ID__n360), .Y(IF_ID__n639) );
  INVx1_ASAP7_75t_R IF_ID___U633 ( .A(IF_ID_inst[17]), .Y(IF_ID__n548) );
  OA21x2_ASAP7_75t_R IF_ID___U634 ( .A1(IF_ID__n525), .A2(IF_ID__n548), .B(IF_ID__n359), .Y(IF_ID__n638) );
  INVx1_ASAP7_75t_R IF_ID___U635 ( .A(IF_ID_inst[18]), .Y(IF_ID__n549) );
  OA21x2_ASAP7_75t_R IF_ID___U636 ( .A1(IF_ID__n525), .A2(IF_ID__n195), .B(IF_ID__n75), .Y(IF_ID__n637) );
  INVx1_ASAP7_75t_R IF_ID___U637 ( .A(IF_ID_inst[19]), .Y(IF_ID__n550) );
  OA21x2_ASAP7_75t_R IF_ID___U638 ( .A1(IF_ID__n526), .A2(IF_ID__n194), .B(IF_ID__n327), .Y(IF_ID__n636) );
  INVx1_ASAP7_75t_R IF_ID___U639 ( .A(IF_ID_inst[20]), .Y(IF_ID__n551) );
  OA21x2_ASAP7_75t_R IF_ID___U640 ( .A1(IF_ID__n526), .A2(IF_ID__n551), .B(IF_ID__n400), .Y(IF_ID__n635) );
  INVx1_ASAP7_75t_R IF_ID___U641 ( .A(IF_ID_inst[21]), .Y(IF_ID__n552) );
  OA21x2_ASAP7_75t_R IF_ID___U642 ( .A1(IF_ID__n527), .A2(IF_ID__n193), .B(IF_ID__n358), .Y(IF_ID__n634) );
  INVx1_ASAP7_75t_R IF_ID___U643 ( .A(IF_ID_inst[22]), .Y(IF_ID__n553) );
  OA21x2_ASAP7_75t_R IF_ID___U644 ( .A1(IF_ID__n527), .A2(IF_ID__n553), .B(IF_ID__n357), .Y(IF_ID__n633) );
  INVx1_ASAP7_75t_R IF_ID___U645 ( .A(IF_ID_inst[23]), .Y(IF_ID__n554) );
  OA21x2_ASAP7_75t_R IF_ID___U646 ( .A1(IF_ID__n2), .A2(IF_ID__n554), .B(IF_ID__IF_ID__n22), .Y(IF_ID__n632) );
  INVx1_ASAP7_75t_R IF_ID___U647 ( .A(IF_ID_inst[24]), .Y(IF_ID__n555) );
  OA21x2_ASAP7_75t_R IF_ID___U648 ( .A1(IF_ID__n527), .A2(IF_ID__n555), .B(IF_ID__n356), .Y(IF_ID__n631) );
  OA21x2_ASAP7_75t_R IF_ID___U649 ( .A1(IF_ID__n119), .A2(IF_ID__n270), .B(IF_ID__n400), .Y(IF_ID__n595) );
  OA21x2_ASAP7_75t_R IF_ID___U650 ( .A1(IF_ID__n1), .A2(IF_ID__n559), .B(IF_ID__n358), .Y(IF_ID__n594) );
  OA21x2_ASAP7_75t_R IF_ID___U651 ( .A1(IF_ID__n528), .A2(IF_ID__n173), .B(IF_ID__n357), .Y(IF_ID__n593) );
  OA21x2_ASAP7_75t_R IF_ID___U652 ( .A1(IF_ID__n529), .A2(IF_ID__n245), .B(IF_ID__n356), .Y(IF_ID__n591) );
  OA21x2_ASAP7_75t_R IF_ID___U653 ( .A1(IF_ID__n12), .A2(IF_ID__n248), .B(IF_ID__n360), .Y(IF_ID__n670) );
  OA21x2_ASAP7_75t_R IF_ID___U654 ( .A1(IF_ID__n1), .A2(IF_ID__n567), .B(IF_ID__n359), .Y(IF_ID__n669) );
  OA21x2_ASAP7_75t_R IF_ID___U655 ( .A1(IF_ID__n527), .A2(IF_ID__n16), .B(IF_ID__n75), .Y(IF_ID__n668) );
  INVx1_ASAP7_75t_R IF_ID___U656 ( .A(IF_ID_rd[0]), .Y(IF_ID__n571) );
  OA21x2_ASAP7_75t_R IF_ID___U657 ( .A1(IF_ID__n12), .A2(IF_ID__n200), .B(IF_ID__n404), .Y(IF_ID__n666) );
  INVx1_ASAP7_75t_R IF_ID___U658 ( .A(IF_ID_rd[1]), .Y(IF_ID__n573) );
  OA21x2_ASAP7_75t_R IF_ID___U659 ( .A1(IF_ID__n527), .A2(IF_ID__n573), .B(IF_ID__n403), .Y(IF_ID__n665) );
  INVx1_ASAP7_75t_R IF_ID___U660 ( .A(IF_ID_rd[2]), .Y(IF_ID__n575) );
  OA21x2_ASAP7_75t_R IF_ID___U661 ( .A1(IF_ID__n527), .A2(IF_ID__n575), .B(IF_ID__n361), .Y(IF_ID__n664) );
  INVx1_ASAP7_75t_R IF_ID___U662 ( .A(IF_ID_rd[3]), .Y(IF_ID__n577) );
  OA21x2_ASAP7_75t_R IF_ID___U663 ( .A1(IF_ID__n12), .A2(IF_ID__IF_ID__n128), .B(IF_ID__n402), .Y(IF_ID__n663) );
  INVx1_ASAP7_75t_R IF_ID___U664 ( .A(IF_ID_rd[4]), .Y(IF_ID__n579) );
  OA21x2_ASAP7_75t_R IF_ID___U665 ( .A1(IF_ID__n530), .A2(IF_ID__n579), .B(IF_ID__n401), .Y(IF_ID__n662) );
  INVx1_ASAP7_75t_R IF_ID___U666 ( .A(IF_ID_opcode[0]), .Y(IF_ID__n581) );
  OA21x2_ASAP7_75t_R IF_ID___U667 ( .A1(IF_ID__n530), .A2(IF_ID__n198), .B(IF_ID__n492), .Y(IF_ID__n661) );
  INVx1_ASAP7_75t_R IF_ID___U668 ( .A(IF_ID_opcode[1]), .Y(IF_ID__n583) );
  OA21x2_ASAP7_75t_R IF_ID___U669 ( .A1(IF_ID__n76), .A2(IF_ID__n237), .B(IF_ID__n407), .Y(IF_ID__n660) );
  OA21x2_ASAP7_75t_R IF_ID___U670 ( .A1(IF_ID__n1), .A2(IF_ID__n586), .B(IF_ID__n363), .Y(IF_ID__n658) );
  OA21x2_ASAP7_75t_R IF_ID___U671 ( .A1(IF_ID__n1), .A2(IF_ID__IF_ID__n143), .B(IF_ID__n405), .Y(IF_ID__n657) );
  OA21x2_ASAP7_75t_R IF_ID___U672 ( .A1(IF_ID__n532), .A2(IF_ID__n589), .B(IF_ID__n376), .Y(IF_ID__n656) );
  OA21x2_ASAP7_75t_R IF_ID___U673 ( .A1(IF_ID__n532), .A2(IF_ID__n235), .B(IF_ID__n362), .Y(IF_ID__n655) );


 
 INVx1_ASAP7_75t_R control___U3 ( .A(control__n32), .Y(control__n9) );
  INVx1_ASAP7_75t_R control___U4 ( .A(control__n4), .Y(control__n34) );
  NAND2x1p5_ASAP7_75t_R control___U5 ( .A(control__n3), .B(control__control__n32), .Y(control__n4) );
  AND5x2_ASAP7_75t_R control___U6 ( .A(opcode[0]), .B(opcode[1]), .C(control__n28), .D(control__n16), .E(
        n20), .Y(control__n32) );
  AND3x2_ASAP7_75t_R control___U7 ( .A(control__n32), .B(opcode[5]), .C(control__n33), .Y(MemWrite) );
  OR2x2_ASAP7_75t_R control___U8 ( .A(opcode[4]), .B(control__n1), .Y(control__n8) );
  NAND2xp33_ASAP7_75t_R control___U9 ( .A(control__n7), .B(control__n28), .Y(control__n1) );
  HB1xp67_ASAP7_75t_R control___U10 ( .A(control__n38), .Y(RegWrite) );
  XNOR2xp5_ASAP7_75t_R control___U11 ( .A(opcode[2]), .B(opcode[3]), .Y(control__n36) );
  HB1xp67_ASAP7_75t_R control___U12 ( .A(control__n24), .Y(control__n20) );
  AOI22xp33_ASAP7_75t_R control___U13 ( .A1(control__n10), .A2(opcode[2]), .B1(control__n11), .B2(control__n12), 
        .Y(control__n24) );
  INVxp67_ASAP7_75t_R control___U14 ( .A(control__n26), .Y(control__n12) );
  HB1xp67_ASAP7_75t_R control___U15 ( .A(control__n25), .Y(control__n26) );
  CKINVDCx20_ASAP7_75t_R control___U16 ( .A(opcode[5]), .Y(control__n3) );
  INVx1_ASAP7_75t_R control___U17 ( .A(control__n8), .Y(control__n5) );
  NAND3xp33_ASAP7_75t_R control___U18 ( .A(opcode[5]), .B(opcode[1]), .C(opcode[0]), .Y(
        n6) );
  INVx1_ASAP7_75t_R control___U19 ( .A(control__n6), .Y(control__n7) );
  INVx1_ASAP7_75t_R control___U20 ( .A(control__n37), .Y(ALUSrc) );
  BUFx2_ASAP7_75t_R control___U21 ( .A(control__n13), .Y(control__n28) );
  INVxp67_ASAP7_75t_R control___U22 ( .A(control__n18), .Y(control__n13) );
  HB1xp67_ASAP7_75t_R control___U23 ( .A(stall), .Y(control__n18) );
  INVxp67_ASAP7_75t_R control___U24 ( .A(opcode[3]), .Y(control__n30) );
  BUFx2_ASAP7_75t_R control___U25 ( .A(control__n21), .Y(control__n25) );
  HB1xp67_ASAP7_75t_R control___U26 ( .A(control__n15), .Y(control__n21) );
  BUFx2_ASAP7_75t_R control___U27 ( .A(control__n17), .Y(control__n16) );
  HB1xp67_ASAP7_75t_R control___U28 ( .A(control__n14), .Y(control__n17) );
  HB1xp67_ASAP7_75t_R control___U29 ( .A(control__n31), .Y(control__n14) );
  XOR2xp5_ASAP7_75t_R control___U30 ( .A(control__n25), .B(opcode[6]), .Y(control__n31) );
  HB1xp67_ASAP7_75t_R control___U31 ( .A(MemtoReg), .Y(MemRead) );
  INVx1_ASAP7_75t_R control___U32 ( .A(control__n23), .Y(control__n11) );
  INVx1_ASAP7_75t_R control___U33 ( .A(control__n30), .Y(control__n10) );
  HB1xp67_ASAP7_75t_R control___U34 ( .A(control__n22), .Y(control__n15) );
  HB1xp67_ASAP7_75t_R control___U35 ( .A(control__n36), .Y(control__n22) );
  OA21x2_ASAP7_75t_R control___U36 ( .A1(opcode[4]), .A2(control__n9), .B(control__n4), .Y(control__n37) );
  BUFx2_ASAP7_75t_R control___U37 ( .A(control__n29), .Y(control__n23) );
  INVx1_ASAP7_75t_R control___U38 ( .A(opcode[6]), .Y(control__n29) );
  AND3x1_ASAP7_75t_R control___U39 ( .A(opcode[6]), .B(control__n5), .C(control__n26), .Y(Branch) );
  INVx3_ASAP7_75t_R control___U40 ( .A(opcode[4]), .Y(control__n33) );
  AND2x2_ASAP7_75t_R control___U41 ( .A(control__n34), .B(control__n33), .Y(MemtoReg) );
  OAI321xp33_ASAP7_75t_R control___U42 ( .A1(control__n8), .A2(control__n16), .A3(control__n20), .B1(control__n9), .B2(control__n33), .C(control__n4), .Y(control__n38) );

  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__25_ ( .D(register__n7631), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[985]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__22_ ( .D(register__n6168), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[982]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__21_ ( .D(register__n7281), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[981]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__20_ ( .D(register__n6514), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[980]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__18_ ( .D(register__n6165), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[978]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__16_ ( .D(register__n6730), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[976]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__8_ ( .D(register__n7282), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[968]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__6_ ( .D(register__n5931), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[966]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__5_ ( .D(register__n7619), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[965]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__4_ ( .D(register__n5708), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[964]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__3_ ( .D(register__n865), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[963]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__2_ ( .D(register__n1485), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[962]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__1_ ( .D(register__n6169), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[961]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__0_ ( .D(register__n947), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[960]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__25_ ( .D(register__n6989), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[953]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__22_ ( .D(register__n878), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[950]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__21_ ( .D(register__n6722), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[949]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__20_ ( .D(register__n9162), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[948]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__16_ ( .D(register__n164), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[944]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__8_ ( .D(register__n757), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[936]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__6_ ( .D(register__n6446), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[934]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__5_ ( .D(register__n1405), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[933]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__4_ ( .D(register__n9163), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[932]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__3_ ( .D(register__n6432), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[931]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__2_ ( .D(register__n7027), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[930]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__1_ ( .D(register__n2174), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[929]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__0_ ( .D(register__n7028), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[928]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__25_ ( .D(register__n4643), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[921]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__22_ ( .D(register__n4383), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[918]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__21_ ( .D(register__n4763), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[917]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__20_ ( .D(register__n735), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[916]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__18_ ( .D(register__n6725), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[914]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__5_ ( .D(register__n4852), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[901]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__4_ ( .D(register__n1156), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[900]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__3_ ( .D(register__n93), .CLK(clk), .SETN(register__n2053), .RESETN(register__n2028), .QN(Reg_data[899]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__0_ ( .D(register__n6731), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[896]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__25_ ( .D(register__n7085), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[857]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__22_ ( .D(register__n805), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[854]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__21_ ( .D(register__n5709), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[853]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__20_ ( .D(register__n5932), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[852]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__18_ ( .D(register__n6170), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[850]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__16_ ( .D(register__n6753), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[848]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__8_ ( .D(register__n7074), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[840]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__6_ ( .D(register__n7075), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[838]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__4_ ( .D(register__net109574), .CLK(clk), 
        .SETN(register__n2053), .RESETN(register__n2028), .QN(Reg_data[836]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__3_ ( .D(register__n6754), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[835]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__2_ ( .D(register__n7076), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[834]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__1_ ( .D(register__n828), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[833]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__0_ ( .D(register__n7029), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[832]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__25_ ( .D(register__n1254), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[825]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__22_ ( .D(register__n7291), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[822]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__21_ ( .D(register__n8646), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[821]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__20_ ( .D(register__n7615), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[820]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__18_ ( .D(register__n8616), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[818]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__16_ ( .D(register__n8596), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[816]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__8_ ( .D(register__n2270), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[808]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__6_ ( .D(register__n1027), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[806]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__5_ ( .D(register__n8617), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[805]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__4_ ( .D(register__n431), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[804]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__2_ ( .D(register__n618), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[802]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__1_ ( .D(register__n788), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[801]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__0_ ( .D(register__n261), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[800]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__25_ ( .D(register__n1051), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[793]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__22_ ( .D(register__n5930), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[790]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__20_ ( .D(register__n476), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[788]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__18_ ( .D(register__n851), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[786]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__16_ ( .D(register__n5234), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[784]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__8_ ( .D(register__n2227), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[776]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__6_ ( .D(register__n1038), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[774]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__5_ ( .D(register__n5379), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[773]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__4_ ( .D(register__n1132), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[772]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__1_ ( .D(register__n1424), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[769]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__0_ ( .D(register__n6755), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[768]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__25_ ( .D(register__n1876), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[761]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__22_ ( .D(register__n5933), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[758]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__21_ ( .D(register__n1077), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[757]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__20_ ( .D(register__n5934), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[756]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__18_ ( .D(register__n4187), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[754]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__16_ ( .D(register__n4277), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[752]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__8_ ( .D(register__n2249), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[744]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__6_ ( .D(register__n4384), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[742]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__5_ ( .D(register__n1367), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[741]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__4_ ( .D(register__n1257), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[740]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__3_ ( .D(register__n5949), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[739]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__2_ ( .D(register__n4589), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[738]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__1_ ( .D(register__n8618), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[737]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__0_ ( .D(register__n1096), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[736]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__25_ ( .D(register__n4764), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[729]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__22_ ( .D(register__n4854), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[726]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__21_ ( .D(register__n1075), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[725]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__20_ ( .D(register__n6171), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[724]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__18_ ( .D(register__n6172), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[722]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__8_ ( .D(register__n2250), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[712]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__6_ ( .D(register__n6173), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[710]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__5_ ( .D(register__n6174), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[709]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__4_ ( .D(register__n6175), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[708]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__3_ ( .D(register__n8648), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[707]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__2_ ( .D(register__n6176), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[706]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__1_ ( .D(register__n5235), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[705]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__0_ ( .D(register__n6177), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[704]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__25_ ( .D(register__n2182), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[697]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__22_ ( .D(register__n610), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[694]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__21_ ( .D(register__n2201), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[693]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__20_ ( .D(register__n2213), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[692]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__18_ ( .D(register__n2196), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[690]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__16_ ( .D(register__n2229), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[688]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__8_ ( .D(register__n2230), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[680]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__6_ ( .D(register__n7893), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[678]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__5_ ( .D(register__n7283), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[677]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__4_ ( .D(register__n7894), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[676]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__3_ ( .D(register__n852), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[675]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__2_ ( .D(register__n7895), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[674]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__1_ ( .D(register__n2219), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[673]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__0_ ( .D(register__n7284), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[672]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__25_ ( .D(register__n1879), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[665]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__22_ ( .D(register__n5547), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[662]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__21_ ( .D(register__n4590), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[661]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__20_ ( .D(register__n4382), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[660]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__18_ ( .D(register__n4275), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[658]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__16_ ( .D(register__n8649), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[656]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__8_ ( .D(register__n4644), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[648]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__6_ ( .D(register__n4765), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[646]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__5_ ( .D(register__n1383), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[645]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__4_ ( .D(register__n325), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[644]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__3_ ( .D(register__n6732), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[643]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__2_ ( .D(register__n9397), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[642]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__1_ ( .D(register__n6726), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[641]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__0_ ( .D(register__n3468), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[640]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__25_ ( .D(register__n296), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[633]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__22_ ( .D(register__n7896), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[630]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__21_ ( .D(register__n7030), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[629]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__20_ ( .D(register__n7897), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[628]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__18_ ( .D(register__n8602), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[626]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__16_ ( .D(register__n7891), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[624]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__8_ ( .D(register__n2271), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[616]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__6_ ( .D(register__n2194), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[614]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__5_ ( .D(register__n7285), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[613]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__4_ ( .D(register__n8673), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[612]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__3_ ( .D(register__n2169), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[611]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__2_ ( .D(register__n1475), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[610]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__1_ ( .D(register__n266), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[609]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__0_ ( .D(register__n2172), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[608]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__25_ ( .D(register__n4855), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[601]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__22_ ( .D(register__n8650), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[598]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__21_ ( .D(register__n602), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[597]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__20_ ( .D(register__n8651), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[596]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__18_ ( .D(register__n4982), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[594]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__16_ ( .D(register__n8652), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[592]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__8_ ( .D(register__n2272), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[584]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__6_ ( .D(register__n1612), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[582]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__5_ ( .D(register__n5236), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[581]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__4_ ( .D(register__n1400), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[580]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__3_ ( .D(register__n6756), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[579]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__2_ ( .D(register__n8653), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[578]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__1_ ( .D(register__n4481), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[577]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__0_ ( .D(register__n5710), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[576]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__25_ ( .D(register__n297), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[569]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__22_ ( .D(register__n3873), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[566]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__21_ ( .D(register__n3911), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[565]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__20_ ( .D(register__n3945), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[564]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__18_ ( .D(register__n3998), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[562]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__16_ ( .D(register__n4048), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[560]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__6_ ( .D(register__n4188), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[550]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__4_ ( .D(register__n4385), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[548]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__3_ ( .D(register__n4486), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[547]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__1_ ( .D(register__n4645), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[545]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__0_ ( .D(register__n4766), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[544]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__25_ ( .D(register__n1362), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[537]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__22_ ( .D(register__n5052), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[534]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__21_ ( .D(register__n283), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[533]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__20_ ( .D(register__n738), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[532]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__18_ ( .D(register__n9403), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[530]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__16_ ( .D(register__n8674), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[528]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__8_ ( .D(register__n2269), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[520]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__6_ ( .D(register__n6200), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[518]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__4_ ( .D(register__n6178), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[516]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__3_ ( .D(register__n5935), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[515]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__2_ ( .D(register__n6179), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[514]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__1_ ( .D(register__n659), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[513]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__0_ ( .D(register__n8592), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[512]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__25_ ( .D(register__n4189), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[473]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__22_ ( .D(register__n5989), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[470]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__21_ ( .D(register__n4156), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[469]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__20_ ( .D(register__n6166), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[468]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__18_ ( .D(register__n6163), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[466]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__16_ ( .D(register__n6180), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[464]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__8_ ( .D(register__n4386), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[456]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__6_ ( .D(register__n4487), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[454]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__4_ ( .D(register__n4591), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[452]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__3_ ( .D(register__n8647), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[451]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__2_ ( .D(register__n9398), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[450]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__0_ ( .D(register__n8603), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[448]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__25_ ( .D(register__n6433), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[441]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__22_ ( .D(register__n8604), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[438]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__21_ ( .D(register__n662), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[437]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__20_ ( .D(register__n2236), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[436]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__18_ ( .D(register__n2200), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[434]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__16_ ( .D(register__n6445), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[432]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__8_ ( .D(register__n2241), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[424]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__6_ ( .D(register__n2237), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[422]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__5_ ( .D(register__n2242), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[421]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__4_ ( .D(register__n4488), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[420]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__3_ ( .D(register__n2240), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[419]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__2_ ( .D(register__n374), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[418]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__1_ ( .D(register__n2191), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[417]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__0_ ( .D(register__n447), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[416]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__25_ ( .D(register__n1870), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[409]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__22_ ( .D(register__n5936), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[406]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__21_ ( .D(register__n661), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[405]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__20_ ( .D(register__n6727), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[404]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__18_ ( .D(register__n9404), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[402]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__16_ ( .D(register__n8675), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[400]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__8_ ( .D(register__n6723), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[392]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__6_ ( .D(register__n1054), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[390]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__5_ ( .D(register__n1425), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[389]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__4_ ( .D(register__n6733), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[388]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__3_ ( .D(register__n9399), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[387]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__2_ ( .D(register__n1423), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[386]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__1_ ( .D(register__n8593), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[385]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__0_ ( .D(register__n445), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[384]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__25_ ( .D(register__n7898), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[377]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__22_ ( .D(register__n1119), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[374]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__21_ ( .D(register__n8605), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[373]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__20_ ( .D(register__n7949), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[372]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__18_ ( .D(register__n3444), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[370]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__16_ ( .D(register__n7892), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[368]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__8_ ( .D(register__n382), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[360]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__6_ ( .D(register__n7950), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[358]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__5_ ( .D(register__n361), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[357]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__4_ ( .D(register__n7031), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[356]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__3_ ( .D(register__n362), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[355]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__2_ ( .D(register__n270), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[354]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__1_ ( .D(register__n384), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[353]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__0_ ( .D(register__n7077), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[352]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__25_ ( .D(register__net122188), .CLK(clk), 
        .SETN(register__n2053), .RESETN(register__n2028), .QN(Reg_data[345]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__22_ ( .D(register__n6201), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[342]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__21_ ( .D(register__n5540), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[341]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__20_ ( .D(register__n8654), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[340]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__18_ ( .D(register__n555), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[338]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__16_ ( .D(register__n8672), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[336]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__8_ ( .D(register__n2226), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[328]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__6_ ( .D(register__n1218), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[326]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__5_ ( .D(register__n7078), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[325]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__4_ ( .D(register__n8671), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[324]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__3_ ( .D(register__n829), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[323]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__2_ ( .D(register__n7084), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[322]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__0_ ( .D(register__n8655), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[320]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__25_ ( .D(register__n3912), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[313]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__22_ ( .D(register__n2263), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[310]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__21_ ( .D(register__n2264), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[309]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__20_ ( .D(register__n2265), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[308]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__18_ ( .D(register__n3872), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[306]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__16_ ( .D(register__n3999), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[304]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__8_ ( .D(register__n4049), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[296]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__5_ ( .D(register__n140), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[293]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__4_ ( .D(register__n4279), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[292]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__3_ ( .D(register__n291), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[291]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__2_ ( .D(register__n6202), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[290]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__1_ ( .D(register__n4387), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[289]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__0_ ( .D(register__n502), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[288]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__25_ ( .D(register__n789), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[281]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__22_ ( .D(register__n8656), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[278]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__21_ ( .D(register__n949), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[277]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__20_ ( .D(register__n6434), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[276]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__18_ ( .D(register__n963), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[274]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__16_ ( .D(register__n1748), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[272]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__8_ ( .D(register__n848), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[264]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__6_ ( .D(register__n4983), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[262]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__5_ ( .D(register__n968), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[261]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__3_ ( .D(register__n6460), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[259]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__2_ ( .D(register__n8657), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[258]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__1_ ( .D(register__n964), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[257]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__0_ ( .D(register__n944), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[256]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__25_ ( .D(register__n7292), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[185]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__22_ ( .D(register__n7286), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[182]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__21_ ( .D(register__n7620), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[181]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__20_ ( .D(register__n1126), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[180]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__18_ ( .D(register__n1263), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[178]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__16_ ( .D(register__n7621), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[176]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__8_ ( .D(register__n1028), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[168]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__6_ ( .D(register__n7287), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[166]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__5_ ( .D(register__n1436), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[165]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__4_ ( .D(register__n1389), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[164]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__3_ ( .D(register__n1125), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[163]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__2_ ( .D(register__n7032), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[162]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__1_ ( .D(register__n7629), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[161]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__0_ ( .D(register__n499), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[160]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__25_ ( .D(register__n1875), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[153]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__22_ ( .D(register__n1487), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[150]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__21_ ( .D(register__n4276), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[149]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__20_ ( .D(register__n4485), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[148]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__18_ ( .D(register__n749), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[146]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__16_ ( .D(register__n4853), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[144]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__8_ ( .D(register__n3406), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[136]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__6_ ( .D(register__n228), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[134]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__4_ ( .D(register__n5937), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[132]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__2_ ( .D(register__n823), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[130]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__1_ ( .D(register__n822), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[129]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__0_ ( .D(register__n511), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[128]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__25_ ( .D(register__n7251), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[121]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__22_ ( .D(register__n6164), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[118]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__21_ ( .D(register__n6681), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[117]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__20_ ( .D(register__n7276), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[116]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__18_ ( .D(register__n7899), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[114]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__16_ ( .D(register__n372), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[112]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__8_ ( .D(register__n7900), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[104]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__5_ ( .D(register__n1686), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[101]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__4_ ( .D(register__n792), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[100]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__3_ ( .D(register__n1689), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[99]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__2_ ( .D(register__n418), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[98]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__1_ ( .D(register__n6682), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[97]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__0_ ( .D(register__n1273), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[96]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__25_ ( .D(register__n7079), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[89]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__22_ ( .D(register__n165), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[86]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__21_ ( .D(register__n7080), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[85]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__20_ ( .D(register__n6203), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[84]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__18_ ( .D(register__n7081), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[82]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__16_ ( .D(register__n138), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[80]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__8_ ( .D(register__n5950), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[72]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__6_ ( .D(register__n7082), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[70]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__5_ ( .D(register__n1055), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[69]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__4_ ( .D(register__n1044), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[68]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__3_ ( .D(register__n6204), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[67]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__2_ ( .D(register__n7083), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[66]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__1_ ( .D(register__n7086), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[65]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__0_ ( .D(register__n1099), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[64]) );
  INVx1_ASAP7_75t_R register___U2084 ( .A(rst), .Y(register__n2053) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__2_ ( .D(register__n7587), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[866]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__0_ ( .D(register__n494), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[864]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__25_ ( .D(register__n2223), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[889]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__22_ ( .D(register__n403), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[886]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__21_ ( .D(register__n5904), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[885]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__1_ ( .D(register__n2238), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[865]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__3_ ( .D(register__n826), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[131]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__20_ ( .D(register__n2209), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[884]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__18_ ( .D(register__n7588), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[882]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__16_ ( .D(register__n386), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[880]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__8_ ( .D(register__n7901), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[872]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__6_ ( .D(register__n7250), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[870]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__5_ ( .D(register__n7252), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[869]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__4_ ( .D(register__n7589), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[868]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__3_ ( .D(register__n7902), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[867]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__16_ ( .D(register__n378), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[16]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__4_ ( .D(register__n5897), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[4]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__2_ ( .D(register__n5948), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[2]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__1_ ( .D(register__n4856), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[1]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__25_ ( .D(register__n5686), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[217]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__22_ ( .D(register__n6181), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[214]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__21_ ( .D(register__n6133), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[213]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__20_ ( .D(register__n4767), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[212]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__18_ ( .D(register__n4984), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[210]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__6_ ( .D(register__n2266), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[198]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__5_ ( .D(register__n5237), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[197]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__4_ ( .D(register__n5380), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[196]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__3_ ( .D(register__n5711), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[195]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__1_ ( .D(register__n5687), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[193]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__0_ ( .D(register__n1176), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[192]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__25_ ( .D(register__n4190), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[25]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__22_ ( .D(register__n4280), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[22]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__20_ ( .D(register__n4388), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[20]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__18_ ( .D(register__n4489), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[18]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__8_ ( .D(register__n4592), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[8]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__6_ ( .D(register__n489), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[6]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__5_ ( .D(register__n4646), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[5]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__8_ ( .D(register__n4857), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[200]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__21_ ( .D(register__n562), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[21]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__2_ ( .D(register__n2294), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[34]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__2_ ( .D(register__n8237), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[226]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__0_ ( .D(register__n6993), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[224]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__25_ ( .D(register__n7590), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[57]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__22_ ( .D(register__n2291), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[54]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__21_ ( .D(register__n8279), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[53]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__25_ ( .D(register__n7033), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[249]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__1_ ( .D(register__n2952), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[225]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__21_ ( .D(register__n7034), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[245]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__16_ ( .D(register__n6182), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[208]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__2_ ( .D(register__n6183), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[194]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__6_ ( .D(register__n449), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[38]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__5_ ( .D(register__n3874), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[37]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__4_ ( .D(register__n1103), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[36]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__3_ ( .D(register__n2740), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[35]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__20_ ( .D(register__n2292), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[244]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__18_ ( .D(register__n7035), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[242]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__8_ ( .D(register__n6126), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[232]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__6_ ( .D(register__n1839), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[230]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__5_ ( .D(register__n13203), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[229]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__4_ ( .D(register__n8238), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[228]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__3_ ( .D(register__n6986), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[227]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__8_ ( .D(register__n7616), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[40]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__16_ ( .D(register__n7036), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[240]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__11_ ( .D(register__n96), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[939]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__11_ ( .D(register__n7617), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[971]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__11_ ( .D(register__n7277), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[811]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__11_ ( .D(register__n351), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[907]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__13_ ( .D(register__n7037), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[813]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__11_ ( .D(register__n6435), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[779]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__11_ ( .D(register__n617), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[107]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__13_ ( .D(register__n131), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[973]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__13_ ( .D(register__n4593), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[301]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__13_ ( .D(register__n6436), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[781]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__11_ ( .D(register__n7038), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[75]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__13_ ( .D(register__n2171), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[621]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__7_ ( .D(register__n1456), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[807]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__7_ ( .D(register__n7278), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[103]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__11_ ( .D(register__n7253), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[619]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__13_ ( .D(register__n5938), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[269]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__11_ ( .D(register__n2293), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[43]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__11_ ( .D(register__n4768), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[11]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__9_ ( .D(register__n9391), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[969]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__31_ ( .D(register__n8595), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[639]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__9_ ( .D(register__n324), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[553]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__7_ ( .D(register__n7622), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[967]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__17_ ( .D(register__n5900), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[881]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__24_ ( .D(register__n8608), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[632]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__13_ ( .D(register__n6437), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[589]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__24_ ( .D(register__n552), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[120]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__7_ ( .D(register__n718), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[775]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__10_ ( .D(register__n426), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[970]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__15_ ( .D(register__n7288), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[687]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__7_ ( .D(register__n6127), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[71]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__7_ ( .D(register__n6734), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[359]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__17_ ( .D(register__n404), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[977]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__11_ ( .D(register__n8658), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[587]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__17_ ( .D(register__n8659), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[625]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__17_ ( .D(register__n5541), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[593]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__28_ ( .D(register__n8678), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[828]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__31_ ( .D(register__n6438), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[991]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__15_ ( .D(register__n1091), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[367]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__13_ ( .D(register__n715), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[45]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__24_ ( .D(register__n6735), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[984]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__30_ ( .D(register__n2208), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[638]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__14_ ( .D(register__n7293), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[622]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__15_ ( .D(register__n7279), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[879]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__9_ ( .D(register__n8609), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[457]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__31_ ( .D(register__n392), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[607]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__13_ ( .D(register__n1688), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[109]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__13_ ( .D(register__n1174), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[77]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__9_ ( .D(register__n390), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[521]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__15_ ( .D(register__n4429), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[975]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__7_ ( .D(register__n2192), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[423]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__17_ ( .D(register__n5216), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[849]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__11_ ( .D(register__n5712), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[523]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__11_ ( .D(register__n4985), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[555]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__24_ ( .D(register__n6736), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[600]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__12_ ( .D(register__n2173), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[620]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__19_ ( .D(register__n173), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[627]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__11_ ( .D(register__n421), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[747]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__11_ ( .D(register__n795), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[875]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__11_ ( .D(register__n3562), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[299]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__11_ ( .D(register__n1109), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[363]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__11_ ( .D(register__n1486), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[395]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__11_ ( .D(register__n2193), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[427]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__11_ ( .D(register__n4647), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[459]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__11_ ( .D(register__n3995), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[651]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__11_ ( .D(register__n4281), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[683]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__11_ ( .D(register__n725), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[715]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__11_ ( .D(register__n1123), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[171]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__11_ ( .D(register__n2284), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[203]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__11_ ( .D(register__n6128), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[235]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__11_ ( .D(register__n6690), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[843]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__11_ ( .D(register__n1008), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[267]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__11_ ( .D(register__n232), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[331]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__11_ ( .D(register__n825), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[139]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__23_ ( .D(register__n7630), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[823]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__27_ ( .D(register__n7039), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[827]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__26_ ( .D(register__n1498), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[634]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__24_ ( .D(register__n6129), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[88]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__30_ ( .D(register__n525), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[62]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__15_ ( .D(register__n8660), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[655]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__30_ ( .D(register__n9392), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[990]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__14_ ( .D(register__n9393), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[974]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__9_ ( .D(register__n5723), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[425]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__28_ ( .D(register__n8680), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[348]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__28_ ( .D(register__n6689), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[988]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__7_ ( .D(register__n7040), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[327]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__31_ ( .D(register__n2211), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[703]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__29_ ( .D(register__n8620), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[189]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__17_ ( .D(register__n251), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[305]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__10_ ( .D(register__n7624), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[810]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__10_ ( .D(register__n6737), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[778]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__19_ ( .D(register__n7654), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[979]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__28_ ( .D(register__n6683), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[796]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__23_ ( .D(register__n357), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[375]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__31_ ( .D(register__n234), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[511]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__15_ ( .D(register__n7041), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[335]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__26_ ( .D(register__n2256), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[890]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__23_ ( .D(register__n7625), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[983]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__13_ ( .D(register__n4046), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[13]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__24_ ( .D(register__n6461), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[312]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__30_ ( .D(register__n8679), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[606]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__14_ ( .D(register__n5637), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[590]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__26_ ( .D(register__n7289), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[986]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__23_ ( .D(register__n8676), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[631]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__23_ ( .D(register__n1573), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[599]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__12_ ( .D(register__n544), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[972]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__15_ ( .D(register__n1395), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[47]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__15_ ( .D(register__n945), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[271]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__7_ ( .D(register__n9183), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[391]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__29_ ( .D(register__n8681), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[317]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__12_ ( .D(register__n6738), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[588]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__19_ ( .D(register__n1252), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[595]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__12_ ( .D(register__n2247), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[876]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__27_ ( .D(register__n4545), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[987]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__13_ ( .D(register__n273), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[365]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__13_ ( .D(register__n306), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[397]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__13_ ( .D(register__n134), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[429]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__13_ ( .D(register__n439), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[461]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__13_ ( .D(register__n7254), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[877]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__13_ ( .D(register__n2243), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[205]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__13_ ( .D(register__n8239), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[237]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__13_ ( .D(register__n1213), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[333]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__13_ ( .D(register__n7026), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[845]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__23_ ( .D(register__n6739), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[791]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_1__29_ ( .D(register__n7325), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[989]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__26_ ( .D(register__n1499), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[602]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__23_ ( .D(register__n7890), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[119]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__13_ ( .D(register__n4769), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[749]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__13_ ( .D(register__n121), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[909]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__13_ ( .D(register__n6684), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[941]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__13_ ( .D(register__n6134), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[525]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__13_ ( .D(register__n487), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[557]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__13_ ( .D(register__n706), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[717]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__28_ ( .D(register__n8682), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[540]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__12_ ( .D(register__n1286), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[460]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__14_ ( .D(register__n4858), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[14]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__30_ ( .D(register__n144), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[382]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__14_ ( .D(register__n853), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[366]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__30_ ( .D(register__n7280), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[126]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__14_ ( .D(register__n423), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[110]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__12_ ( .D(register__n2295), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[44]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__12_ ( .D(register__n7042), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[236]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__13_ ( .D(register__n723), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[141]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__13_ ( .D(register__n2248), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[173]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__13_ ( .D(register__n4047), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[653]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__13_ ( .D(register__n6396), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[685]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__9_ ( .D(register__n8663), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[393]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__28_ ( .D(register__n7952), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[380]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__28_ ( .D(register__n8281), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[252]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__31_ ( .D(register__n238), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[671]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__29_ ( .D(register__n1497), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[157]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__7_ ( .D(register__n2170), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[615]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__7_ ( .D(register__n5939), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[583]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__17_ ( .D(register__n6439), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[273]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__25_ ( .D(register__n3639), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[505]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__12_ ( .D(register__n3753), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[556]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__19_ ( .D(register__n409), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[403]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__7_ ( .D(register__n2296), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[39]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__7_ ( .D(register__n2260), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[199]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__7_ ( .D(register__n6399), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[231]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__7_ ( .D(register__n5542), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[263]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__10_ ( .D(register__n7903), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[618]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__23_ ( .D(register__n8610), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[343]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__31_ ( .D(register__n6190), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[479]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__27_ ( .D(register__n6184), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[539]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__23_ ( .D(register__n3997), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[439]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__26_ ( .D(register__n6740), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[858]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__24_ ( .D(register__n8664), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[280]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__16_ ( .D(register__n143), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[496]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__22_ ( .D(register__n604), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[502]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__20_ ( .D(register__n4594), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[500]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__18_ ( .D(register__n356), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[498]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__13_ ( .D(register__n510), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[493]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__12_ ( .D(register__n4859), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[492]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__11_ ( .D(register__n163), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[491]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__9_ ( .D(register__n4986), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[489]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__8_ ( .D(register__n591), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[488]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__6_ ( .D(register__n5053), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[486]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__5_ ( .D(register__n7326), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[485]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__4_ ( .D(register__n3082), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[484]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__2_ ( .D(register__n5381), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[482]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__0_ ( .D(register__n3081), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[480]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__26_ ( .D(register__n4648), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[314]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__26_ ( .D(register__n8280), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[250]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__21_ ( .D(register__n607), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[501]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__1_ ( .D(register__n3050), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[481]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__12_ ( .D(register__n4770), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[300]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__15_ ( .D(register__n4860), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[303]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__27_ ( .D(register__n6741), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[411]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__29_ ( .D(register__n1227), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[285]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__9_ ( .D(register__n619), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[617]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__9_ ( .D(register__n2231), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[681]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__29_ ( .D(register__n7905), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[125]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__29_ ( .D(register__n8683), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[253]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__17_ ( .D(register__n2273), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[817]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__31_ ( .D(register__n6135), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[543]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__9_ ( .D(register__n8611), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[809]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__9_ ( .D(register__n379), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[873]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__9_ ( .D(register__n3663), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[137]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__9_ ( .D(register__n7626), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[169]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__9_ ( .D(register__n777), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[777]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__9_ ( .D(register__n6742), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[841]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__31_ ( .D(register__n148), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[575]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__28_ ( .D(register__n7632), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[572]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__17_ ( .D(register__n444), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[113]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__17_ ( .D(register__n6185), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[81]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__24_ ( .D(register__n5906), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[536]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__24_ ( .D(register__n737), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[568]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__12_ ( .D(register__n9400), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[204]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__12_ ( .D(register__n2165), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[12]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__30_ ( .D(register__n7051), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[94]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__30_ ( .D(register__n130), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[350]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__14_ ( .D(register__n8665), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[334]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__31_ ( .D(register__n5218), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[415]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__31_ ( .D(register__n4979), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[447]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__28_ ( .D(register__n7953), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[220]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__24_ ( .D(register__n8612), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[376]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__24_ ( .D(register__n6728), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[408]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__24_ ( .D(register__n160), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[56]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__24_ ( .D(register__n2168), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[216]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__24_ ( .D(register__n8240), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[248]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__24_ ( .D(register__n4987), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[24]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__24_ ( .D(register__net119141), .CLK(clk), 
        .SETN(register__n2053), .RESETN(register__n2028), .QN(Reg_data[344]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__24_ ( .D(register__n1752), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[440]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__15_ ( .D(register__n2128), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[751]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__15_ ( .D(register__n6994), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[815]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__15_ ( .D(register__n4981), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[911]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__15_ ( .D(register__n1406), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[943]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__15_ ( .D(register__n824), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[143]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__15_ ( .D(register__n6685), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[175]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__15_ ( .D(register__n6167), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[527]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__15_ ( .D(register__n246), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[559]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__15_ ( .D(register__n4482), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[719]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__15_ ( .D(register__n4642), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[591]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__15_ ( .D(register__n363), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[783]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__15_ ( .D(register__n7043), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[623]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__12_ ( .D(register__n1293), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[524]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__15_ ( .D(register__n5713), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[207]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__15_ ( .D(register__n6401), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[239]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__15_ ( .D(register__n365), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[399]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__15_ ( .D(register__n1023), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[431]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__15_ ( .D(register__n5714), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[495]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__15_ ( .D(register__n1020), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[111]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__15_ ( .D(register__n1404), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[79]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__19_ ( .D(register__n2164), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[19]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__10_ ( .D(register__n2934), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[586]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__15_ ( .D(register__n4861), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[463]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__19_ ( .D(register__n1855), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[435]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__3_ ( .D(register__n5940), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[483]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__23_ ( .D(register__n354), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[407]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__27_ ( .D(register__n5239), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[571]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__26_ ( .D(register__n9401), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[218]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__26_ ( .D(register__n6440), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[282]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__12_ ( .D(register__n8668), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[268]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__7_ ( .D(register__n5901), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[743]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__7_ ( .D(register__n7591), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[871]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__7_ ( .D(register__n5370), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[903]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__7_ ( .D(register__n9164), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[935]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__7_ ( .D(register__n501), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[135]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__7_ ( .D(register__n1241), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[167]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__7_ ( .D(register__n5941), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[519]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__7_ ( .D(register__n5382), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[551]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__7_ ( .D(register__n5054), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[647]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__7_ ( .D(register__n6990), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[679]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__7_ ( .D(register__n5219), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[711]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__7_ ( .D(register__net111717), .CLK(clk), 
        .SETN(register__n2053), .RESETN(register__n2028), .QN(Reg_data[839]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__28_ ( .D(register__n1064), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[636]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__28_ ( .D(register__n1062), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[604]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__27_ ( .D(register__n2239), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[443]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__7_ ( .D(register__n4183), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[455]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__7_ ( .D(register__n3592), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[487]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__9_ ( .D(register__n8669), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[585]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__9_ ( .D(register__n8670), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[649]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__30_ ( .D(register__n7951), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[318]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__14_ ( .D(register__n3836), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[302]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__30_ ( .D(register__n166), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[222]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__14_ ( .D(register__n870), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[206]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__30_ ( .D(register__n6997), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[254]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__14_ ( .D(register__n7044), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[238]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__30_ ( .D(register__n962), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[286]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__14_ ( .D(register__n5715), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[270]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__29_ ( .D(register__n9402), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[221]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__29_ ( .D(register__n803), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[93]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__30_ ( .D(register__n8597), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[574]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__30_ ( .D(register__n2176), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[766]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__14_ ( .D(register__n609), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[750]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__30_ ( .D(register__n8677), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[830]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__14_ ( .D(register__n2084), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[814]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__30_ ( .D(register__n7255), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[894]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__14_ ( .D(register__n5905), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[878]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__30_ ( .D(register__n9394), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[926]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__14_ ( .D(register__n886), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[910]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__30_ ( .D(register__n7025), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[958]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__14_ ( .D(register__n873), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[942]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__30_ ( .D(register__n850), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[158]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__14_ ( .D(register__n4588), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[142]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__30_ ( .D(register__n7256), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[190]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__14_ ( .D(register__n1056), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[174]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__30_ ( .D(register__n8621), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[542]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__14_ ( .D(register__n5907), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[526]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__14_ ( .D(register__n7049), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[558]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__30_ ( .D(register__n135), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[670]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__14_ ( .D(register__n5240), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[654]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__30_ ( .D(register__n2183), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[702]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__14_ ( .D(register__n7871), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[686]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__30_ ( .D(register__n8582), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[734]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__14_ ( .D(register__n542), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[718]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__30_ ( .D(register__n7294), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[798]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__14_ ( .D(register__n854), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[782]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__30_ ( .D(register__n624), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[862]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__14_ ( .D(register__n7048), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[846]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__17_ ( .D(register__n2297), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[785]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__10_ ( .D(register__n5055), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[746]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__10_ ( .D(register__n614), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[874]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__10_ ( .D(register__n1253), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[906]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__10_ ( .D(register__n1250), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[938]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__10_ ( .D(register__n1121), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[170]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__10_ ( .D(register__n6136), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[522]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__10_ ( .D(register__n6743), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[650]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__10_ ( .D(register__n2181), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[682]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__10_ ( .D(register__n5220), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[714]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__10_ ( .D(register__n7045), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[842]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__10_ ( .D(register__n5543), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[554]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__28_ ( .D(register__n95), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[316]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__28_ ( .D(register__n6691), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[412]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__28_ ( .D(register__n5369), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[476]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__28_ ( .D(register__n8684), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[508]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__28_ ( .D(register__n2287), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[60]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__28_ ( .D(register__n6696), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[124]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__28_ ( .D(register__n4988), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[28]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__28_ ( .D(register__n1221), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[92]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__28_ ( .D(register__n948), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[284]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__28_ ( .D(register__n8583), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[444]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__12_ ( .D(register__n5241), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[748]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__12_ ( .D(register__n7627), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[812]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__12_ ( .D(register__n595), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[908]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__12_ ( .D(register__n9165), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[940]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__12_ ( .D(register__n1078), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[140]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__12_ ( .D(register__n7628), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[172]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__12_ ( .D(register__n5383), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[652]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__12_ ( .D(register__n2204), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[684]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__12_ ( .D(register__n4585), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[716]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__12_ ( .D(register__n5716), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[780]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__19_ ( .D(register__n4989), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[307]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__19_ ( .D(register__n9395), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[371]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__19_ ( .D(register__n5371), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[467]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__19_ ( .D(register__n1223), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[755]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__19_ ( .D(register__n6995), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[819]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__19_ ( .D(register__n7873), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[883]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__19_ ( .D(register__n508), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[915]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__19_ ( .D(register__n2175), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[947]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__19_ ( .D(register__n6400), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[115]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__19_ ( .D(register__n5942), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[211]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__19_ ( .D(register__n8241), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[243]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__19_ ( .D(register__n3404), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[147]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__19_ ( .D(register__n1157), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[179]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__19_ ( .D(register__n5544), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[531]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__19_ ( .D(register__n4184), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[659]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__19_ ( .D(register__n5221), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[723]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__19_ ( .D(register__n6186), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[83]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__19_ ( .D(register__n5943), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[275]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__19_ ( .D(register__n5944), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[339]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__19_ ( .D(register__n6442), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[851]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__19_ ( .D(register__n391), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[499]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__19_ ( .D(register__n5717), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[563]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__19_ ( .D(register__n2198), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[691]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__10_ ( .D(register__n3640), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[298]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__10_ ( .D(register__n352), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[362]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__10_ ( .D(register__n6692), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[394]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__10_ ( .D(register__n4990), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[458]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__10_ ( .D(register__n3870), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[490]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__10_ ( .D(register__n1310), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[42]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__10_ ( .D(register__n4191), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[106]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__10_ ( .D(register__n2283), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[202]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__10_ ( .D(register__n6402), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[234]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__10_ ( .D(register__n5056), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[10]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__10_ ( .D(register__n5384), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[74]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__10_ ( .D(register__n6403), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[266]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__10_ ( .D(register__n5902), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[330]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__10_ ( .D(register__n2221), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[426]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__23_ ( .D(register__n4584), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[759]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__23_ ( .D(register__n7248), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[887]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__23_ ( .D(register__n551), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[919]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__23_ ( .D(register__n1305), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[951]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__23_ ( .D(register__n819), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[151]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__23_ ( .D(register__n1392), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[183]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__23_ ( .D(register__n6137), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[535]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__23_ ( .D(register__n5945), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[567]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__23_ ( .D(register__n4126), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[663]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__23_ ( .D(register__n2184), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[695]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__23_ ( .D(register__n5385), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[727]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__23_ ( .D(register__n1173), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[855]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__27_ ( .D(register__n8594), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[763]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__27_ ( .D(register__n2255), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[891]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__27_ ( .D(register__n322), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[923]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__27_ ( .D(register__n313), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[955]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__27_ ( .D(register__n4186), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[155]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__27_ ( .D(register__n299), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[187]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__27_ ( .D(register__n295), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[635]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__27_ ( .D(register__n310), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[667]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__27_ ( .D(register__n2178), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[699]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__27_ ( .D(register__n4762), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[603]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__27_ ( .D(register__net109491), .CLK(clk), 
        .SETN(register__n2053), .RESETN(register__n2028), .QN(Reg_data[859]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__23_ ( .D(register__n5057), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[311]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__23_ ( .D(register__n5058), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[471]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__23_ ( .D(register__n4381), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[503]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__23_ ( .D(register__n1072), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[55]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__23_ ( .D(register__n5707), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[215]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__23_ ( .D(register__n5242), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[23]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__23_ ( .D(register__n1009), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[279]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__27_ ( .D(register__n8598), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[731]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__9_ ( .D(register__n8613), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[361]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__9_ ( .D(register__n6130), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[41]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__9_ ( .D(register__n6694), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[105]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__9_ ( .D(register__n2133), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[201]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__9_ ( .D(register__n776), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[233]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__9_ ( .D(register__n5386), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[9]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__9_ ( .D(register__n6187), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[265]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__9_ ( .D(register__n5946), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[329]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__26_ ( .D(register__n5908), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[762]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__26_ ( .D(register__n7249), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[826]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__26_ ( .D(register__n755), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[922]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__26_ ( .D(register__n9166), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[954]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__26_ ( .D(register__n3834), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[154]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__26_ ( .D(register__n6686), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[186]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__26_ ( .D(register__n529), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[538]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__26_ ( .D(register__n6188), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[570]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__26_ ( .D(register__n6744), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[666]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__26_ ( .D(register__n2177), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[698]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__26_ ( .D(register__n6131), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[730]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__26_ ( .D(register__n6189), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[794]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__31_ ( .D(register__n240), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[767]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__31_ ( .D(register__n7618), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[831]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__31_ ( .D(register__n5372), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[927]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__31_ ( .D(register__n9184), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[959]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__31_ ( .D(register__n654), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[159]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__31_ ( .D(register__n1396), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[191]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__31_ ( .D(register__n1086), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[735]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__31_ ( .D(register__n6996), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[799]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__31_ ( .D(register__n1152), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[863]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__9_ ( .D(register__n5545), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[745]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__9_ ( .D(register__n1560), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[905]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__9_ ( .D(register__n97), .CLK(clk), .SETN(register__n2053), .RESETN(register__n2028), .QN(Reg_data[937]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__9_ ( .D(register__n6138), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[713]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__26_ ( .D(register__n383), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[378]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__26_ ( .D(register__n5909), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[410]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__26_ ( .D(register__n5243), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[442]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__26_ ( .D(register__n5244), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[474]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__26_ ( .D(register__n3079), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[506]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__26_ ( .D(register__n1016), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[122]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__26_ ( .D(register__n1018), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[90]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__26_ ( .D(register__n4973), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[346]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__12_ ( .D(register__n8614), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[364]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__12_ ( .D(register__n5911), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[396]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__12_ ( .D(register__n92), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[428]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__12_ ( .D(register__n1015), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[108]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__12_ ( .D(register__n5718), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[76]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__12_ ( .D(register__n7046), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[332]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__17_ ( .D(register__n408), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[945]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__17_ ( .D(register__n1401), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[177]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__17_ ( .D(register__n5719), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[753]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__17_ ( .D(register__n6729), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[913]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__17_ ( .D(register__n5539), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[145]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__17_ ( .D(register__n5910), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[529]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__17_ ( .D(register__n6443), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[561]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__17_ ( .D(register__n6688), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[657]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__17_ ( .D(register__n2179), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[689]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__17_ ( .D(register__n6132), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[721]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__17_ ( .D(register__n8555), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[369]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__17_ ( .D(register__n5373), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[401]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__17_ ( .D(register__n255), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[465]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__17_ ( .D(register__n484), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[497]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__17_ ( .D(register__n6444), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[209]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__17_ ( .D(register__n8242), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[241]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__17_ ( .D(register__n1017), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[337]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__24_ ( .D(register__n937), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[760]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__24_ ( .D(register__n8615), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[824]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__24_ ( .D(register__n2210), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[888]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__24_ ( .D(register__n5947), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[920]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__24_ ( .D(register__n9167), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[952]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__24_ ( .D(register__n3871), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[152]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__24_ ( .D(register__n6991), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[184]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__24_ ( .D(register__n6687), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[664]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__24_ ( .D(register__n2180), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[696]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__24_ ( .D(register__n943), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[728]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__24_ ( .D(register__n736), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[792]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__24_ ( .D(register__n938), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[856]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__27_ ( .D(register__n5387), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[315]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__27_ ( .D(register__n5388), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[475]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__27_ ( .D(register__n7290), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[123]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__27_ ( .D(register__n282), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[251]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__27_ ( .D(register__n7047), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[91]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__27_ ( .D(register__n950), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[283]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__27_ ( .D(register__net109782), .CLK(clk), 
        .SETN(register__n2053), .RESETN(register__n2028), .QN(Reg_data[347]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__27_ ( .D(register__n330), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[379]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__27_ ( .D(register__n225), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[219]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__31_ ( .D(register__n8556), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[319]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__31_ ( .D(register__n6693), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[383]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__31_ ( .D(register__n7872), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[127]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_25__31_ ( .D(register__n4586), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[223]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__31_ ( .D(register__n8243), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[255]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__31_ ( .D(register__n4846), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[31]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__31_ ( .D(register__n132), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[95]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__31_ ( .D(register__n967), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[287]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__31_ ( .D(register__n8599), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[351]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__29_ ( .D(register__n2289), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[61]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_20__29_ ( .D(register__n8685), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[381]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__29_ ( .D(register__n1871), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[413]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__29_ ( .D(register__n961), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[445]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__29_ ( .D(register__n1236), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[477]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__29_ ( .D(register__n1235), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[509]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__29_ ( .D(register__n5903), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[29]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__29_ ( .D(register__n1574), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[349]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__29_ ( .D(register__n7655), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[829]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__29_ ( .D(register__n847), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[765]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__29_ ( .D(register__n2218), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[893]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__29_ ( .D(register__n7904), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[925]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__29_ ( .D(register__n6695), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[957]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__29_ ( .D(register__n2267), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[541]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__29_ ( .D(register__n8622), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[573]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_12__29_ ( .D(register__n6992), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[637]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__29_ ( .D(register__n8623), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[669]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__29_ ( .D(register__n1231), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[701]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__29_ ( .D(register__n5222), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[733]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_13__29_ ( .D(register__n1609), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[605]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__29_ ( .D(register__n332), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[797]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__29_ ( .D(register__n5217), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[861]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_8__28_ ( .D(register__n8624), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[764]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__28_ ( .D(register__n161), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[892]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__28_ ( .D(register__n5374), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[924]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__28_ ( .D(register__n9185), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[956]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__28_ ( .D(register__n613), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[156]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_26__28_ ( .D(register__n298), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[188]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_11__28_ ( .D(register__n1065), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[668]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_10__28_ ( .D(register__n563), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[700]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__28_ ( .D(register__n170), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[860]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__28_ ( .D(register__n8625), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[732]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__30_ ( .D(register__n440), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[446]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__30_ ( .D(register__n438), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[414]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_19__14_ ( .D(register__n2257), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[398]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__30_ ( .D(register__n1079), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[478]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__14_ ( .D(register__n5546), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[462]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__30_ ( .D(register__n371), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[510]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__14_ ( .D(register__n3942), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[494]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__6_ ( .D(register__n2085), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[902]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__27_ ( .D(register__n2074), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[27]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__17_ ( .D(register__n2073), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[17]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__3_ ( .D(register__n2072), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[3]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_2__18_ ( .D(register__n9388), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[946]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__14_ ( .D(register__n2071), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[430]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_18__17_ ( .D(register__n2070), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[433]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__15_ ( .D(register__n2069), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[15]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__6_ ( .D(register__n2068), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[294]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__20_ ( .D(register__n2067), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[52]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__19_ ( .D(register__n2066), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[51]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__18_ ( .D(register__n2065), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[50]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__17_ ( .D(register__n2064), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[49]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__1_ ( .D(register__n2063), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[33]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__7_ ( .D(register__n2062), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[7]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__7_ ( .D(register__n2061), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[295]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__10_ ( .D(register__n2060), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[138]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__2_ ( .D(register__n2059), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[546]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__0_ ( .D(register__n167), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[0]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__27_ ( .D(register__n2058), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[795]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__1_ ( .D(register__n289), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[897]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__0_ ( .D(register__n2057), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[32]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__2_ ( .D(register__n2056), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[898]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_22__9_ ( .D(register__n2055), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[297]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__12_ ( .D(register__n2054), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[844]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_4__31_ ( .D(register__n2232), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[895]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__31_ ( .D(register__n2290), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[63]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__27_ ( .D(register__n936), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[59]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_28__6_ ( .D(register__n395), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[102]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__2_ ( .D(register__n2052), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[770]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__5_ ( .D(register__net111561), .CLK(clk), 
        .SETN(register__n2053), .RESETN(register__n2028), .QN(Reg_data[837]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__16_ ( .D(register__n2288), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[48]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__8_ ( .D(register__n2051), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[552]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_23__4_ ( .D(register__n2050), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[260]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__26_ ( .D(register__n2049), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[26]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_9__16_ ( .D(register__n2048), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[720]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__14_ ( .D(register__n2047), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[46]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__21_ ( .D(register__n2046), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[789]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_6__3_ ( .D(register__n2045), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[803]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_30__26_ ( .D(register__n2044), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[58]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__23_ ( .D(register__n2043), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[87]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__14_ ( .D(register__n512), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[78]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__5_ ( .D(register__n2042), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[453]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_14__5_ ( .D(register__n2041), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[549]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__16_ ( .D(register__n2040), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[912]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_29__9_ ( .D(register__n2039), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[73]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__1_ ( .D(register__n2038), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[449]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__3_ ( .D(register__n2037), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[771]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_21__1_ ( .D(register__n2036), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[321]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_31__30_ ( .D(register__n2035), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[30]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_7__19_ ( .D(register__n2034), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[787]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_27__5_ ( .D(register__n2033), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[133]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__24_ ( .D(register__n2032), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[504]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_15__5_ ( .D(register__n2268), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[517]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_17__24_ ( .D(register__n2031), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[472]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_16__27_ ( .D(register__n314), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[507]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_5__15_ ( .D(register__n2030), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[847]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_3__8_ ( .D(register__n2079), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[904]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__23_ ( .D(register__n2029), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[247]) );
  DFFASRHQNx1_ASAP7_75t_R register___Reg_data_reg_24__22_ ( .D(register__n2027), .CLK(clk), .SETN(
        n2053), .RESETN(register__n2028), .QN(Reg_data[246]) );
  TIEHIx1_ASAP7_75t_R register___U2 ( .H(register__n2028) );
  INVxp67_ASAP7_75t_R register___U3 ( .A(register__n11116), .Y(register__n5928) );
  INVxp67_ASAP7_75t_R register___U4 ( .A(register__n10854), .Y(register__n5913) );
  INVxp67_ASAP7_75t_R register___U5 ( .A(register__n10610), .Y(register__n7909) );
  AOI21xp5_ASAP7_75t_R register___U6 ( .A1(register__n281), .A2(register__net89993), .B(register__n2343), .Y(register__n2364) );
  OR2x4_ASAP7_75t_R register___U7 ( .A(register__n1104), .B(register__n14), .Y(register__n327) );
  INVx4_ASAP7_75t_R register___U8 ( .A(IF_ID_rs1[3]), .Y(register__n11150) );
  CKINVDCx10_ASAP7_75t_R register___U9 ( .A(register__C6422_net59546), .Y(register__n2002) );
  AND2x6_ASAP7_75t_R register___U10 ( .A(IF_ID_rs1[4]), .B(register__n56), .Y(register__n1226) );
  INVx1_ASAP7_75t_R register___U11 ( .A(register__n1863), .Y(register__n1864) );
  BUFx4f_ASAP7_75t_R register___U12 ( .A(register__n885), .Y(register__n1) );
  INVx1_ASAP7_75t_R register___U13 ( .A(register__n1247), .Y(register__n2) );
  INVx2_ASAP7_75t_R register___U14 ( .A(register__net120788), .Y(register__n1247) );
  AND2x6_ASAP7_75t_R register___U15 ( .A(register__n13), .B(register__n11149), .Y(register__n3) );
  AND2x6_ASAP7_75t_R register___U16 ( .A(register__n565), .B(register__n8752), .Y(register__n11149) );
  AND2x2_ASAP7_75t_R register___U17 ( .A(register__net126601), .B(register__net89045), .Y(register__n4) );
  NOR2xp67_ASAP7_75t_R register___U18 ( .A(register__n4), .B(register__n2669), .Y(register__n2671) );
  BUFx6f_ASAP7_75t_R register___U19 ( .A(register__net89046), .Y(register__net89045) );
  INVx6_ASAP7_75t_R register___U20 ( .A(register__net117657), .Y(register__n1398) );
  AO22x1_ASAP7_75t_R register___U21 ( .A1(register__n50), .A2(register__n2235), .B1(register__n1851), .B2(register__n2234), .Y(
        read_reg_data_1[26]) );
  INVx1_ASAP7_75t_R register___U22 ( .A(register__n5278), .Y(register__n6) );
  BUFx4f_ASAP7_75t_R register___U23 ( .A(register__n4933), .Y(register__n4932) );
  NOR2x1_ASAP7_75t_R register___U24 ( .A(register__n3104), .B(register__n3103), .Y(register__n35) );
  OAI22xp33_ASAP7_75t_R register___U25 ( .A1(register__n53), .A2(register__n8644), .B1(register__net61369), .B2(
        net64696), .Y(read_reg_data_1[7]) );
  INVx3_ASAP7_75t_R register___U26 ( .A(register__net131160), .Y(register__n388) );
  INVxp67_ASAP7_75t_R register___U27 ( .A(register__n5458), .Y(register__n7) );
  INVx6_ASAP7_75t_R register___U28 ( .A(register__net126601), .Y(register__net109643) );
  AOI22xp5_ASAP7_75t_R register___U29 ( .A1(register__n8753), .A2(register__net146144), .B1(register__n10229), .B2(
        net126601), .Y(register__n705) );
  NOR2xp67_ASAP7_75t_R register___U30 ( .A(register__n1117), .B(register__net109872), .Y(register__n253) );
  INVx4_ASAP7_75t_R register___U31 ( .A(register__n1996), .Y(register__n1117) );
  OR2x2_ASAP7_75t_R register___U32 ( .A(register__C6422_net59729), .B(register__n2002), .Y(register__n561) );
  INVx1_ASAP7_75t_R register___U33 ( .A(register__n5459), .Y(register__n8) );
  NOR2x1_ASAP7_75t_R register___U34 ( .A(register__n2373), .B(register__n2374), .Y(register__n2395) );
  INVx1_ASAP7_75t_R register___U35 ( .A(register__n10701), .Y(register__n9) );
  AND2x2_ASAP7_75t_R register___U36 ( .A(register__n1996), .B(register__C6423_net60596), .Y(register__n941) );
  CKINVDCx9p33_ASAP7_75t_R register___U37 ( .A(register__n1996), .Y(register__n1997) );
  NAND2xp33_ASAP7_75t_R register___U38 ( .A(register__n2766), .B(register__n8747), .Y(register__n11) );
  OR2x2_ASAP7_75t_R register___U39 ( .A(register__n1330), .B(register__n237), .Y(register__n10) );
  AO22x1_ASAP7_75t_R register___U40 ( .A1(register__n52), .A2(register__n11), .B1(register__n1851), .B2(register__net62656), .Y(
        read_reg_data_1[31]) );
  INVx2_ASAP7_75t_R register___U41 ( .A(register__net62684), .Y(register__net62656) );
  INVx1_ASAP7_75t_R register___U42 ( .A(register__n5454), .Y(register__n12) );
  INVx3_ASAP7_75t_R register___U43 ( .A(register__n1577), .Y(register__n1578) );
  BUFx6f_ASAP7_75t_R register___U44 ( .A(register__n381), .Y(register__n233) );
  BUFx12f_ASAP7_75t_R register___U45 ( .A(register__n387), .Y(register__net131160) );
  OAI22xp33_ASAP7_75t_R register___U46 ( .A1(register__n54), .A2(register__n7024), .B1(register__net61369), .B2(
        net141997), .Y(read_reg_data_1[23]) );
  INVx2_ASAP7_75t_R register___U47 ( .A(register__n507), .Y(register__n1909) );
  INVx2_ASAP7_75t_R register___U48 ( .A(register__n5032), .Y(register__n7605) );
  AOI21xp33_ASAP7_75t_R register___U49 ( .A1(register__n39), .A2(register__net90253), .B(register__n2666), .Y(register__n2668) );
  NAND2xp67_ASAP7_75t_R register___U50 ( .A(register__n2769), .B(register__n779), .Y(register__n2235) );
  BUFx3_ASAP7_75t_R register___U51 ( .A(register__n4922), .Y(register__n4921) );
  NAND2xp5_ASAP7_75t_R register___U52 ( .A(register__n2746), .B(register__n10818), .Y(register__n226) );
  BUFx12f_ASAP7_75t_R register___U53 ( .A(register__n437), .Y(register__n13) );
  AND2x4_ASAP7_75t_R register___U54 ( .A(IF_ID_rs1[4]), .B(register__n11150), .Y(register__n437) );
  INVxp67_ASAP7_75t_R register___U55 ( .A(register__n437), .Y(register__n222) );
  NOR2xp67_ASAP7_75t_R register___U56 ( .A(register__n2647), .B(register__n2646), .Y(register__n2670) );
  NAND2xp5_ASAP7_75t_R register___U57 ( .A(register__register__n11153), .B(register__n1), .Y(register__register__n14) );
  INVx2_ASAP7_75t_R register___U58 ( .A(IF_ID_rs1[4]), .Y(register__n11153) );
  OR2x2_ASAP7_75t_R register___U59 ( .A(register__net117656), .B(register__n2331), .Y(register__n15) );
  CKINVDCx8_ASAP7_75t_R register___U60 ( .A(register__n817), .Y(register__n1996) );
  INVx6_ASAP7_75t_R register___U61 ( .A(register__C6422_net59540), .Y(register__n802) );
  INVx4_ASAP7_75t_R register___U62 ( .A(register__C6422_net59540), .Y(register__n801) );
  OR2x2_ASAP7_75t_R register___U63 ( .A(register__C6422_net59726), .B(register__n800), .Y(register__n16) );
  OR2x2_ASAP7_75t_R register___U64 ( .A(register__n66), .B(register__n2637), .Y(register__n17) );
  BUFx4f_ASAP7_75t_R register___U65 ( .A(register__net139537), .Y(register__C6422_net70296) );
  CKINVDCx8_ASAP7_75t_R register___U66 ( .A(register__n327), .Y(register__net123857) );
  INVx6_ASAP7_75t_R register___U67 ( .A(register__n381), .Y(register__n1577) );
  INVx2_ASAP7_75t_R register___U68 ( .A(register__n1577), .Y(register__n1579) );
  INVx3_ASAP7_75t_R register___U69 ( .A(register__C6422_net70602), .Y(register__n1420) );
  OR2x2_ASAP7_75t_R register___U70 ( .A(register__net64864), .B(register__net61369), .Y(register__n18) );
  OR2x2_ASAP7_75t_R register___U71 ( .A(register__net61369), .B(register__n12249), .Y(register__n19) );
  INVx4_ASAP7_75t_R register___U72 ( .A(register__n55), .Y(register__n48) );
  CKINVDCx5p33_ASAP7_75t_R register___U73 ( .A(register__n52), .Y(register__n53) );
  INVx4_ASAP7_75t_R register___U74 ( .A(register__n50), .Y(register__n54) );
  INVx3_ASAP7_75t_R register___U75 ( .A(register__n48), .Y(register__n52) );
  INVxp67_ASAP7_75t_R register___U76 ( .A(register__n48), .Y(register__n51) );
  INVx2_ASAP7_75t_R register___U77 ( .A(register__n48), .Y(register__n50) );
  XNOR2x2_ASAP7_75t_R register___U78 ( .A(register__n11847), .B(register__n4264), .Y(register__n12515) );
  INVx2_ASAP7_75t_R register___U79 ( .A(register__n368), .Y(register__n369) );
  BUFx4f_ASAP7_75t_R register___U80 ( .A(register__C6422_net60443), .Y(register__C6422_net70678) );
  INVx4_ASAP7_75t_R register___U81 ( .A(register__net120912), .Y(register__n1336) );
  BUFx2_ASAP7_75t_R register___U82 ( .A(register__n11028), .Y(register__n5957) );
  BUFx6f_ASAP7_75t_R register___U83 ( .A(register__net120912), .Y(register__n326) );
  INVx3_ASAP7_75t_R register___U84 ( .A(register__C6422_net59538), .Y(register__n419) );
  BUFx2_ASAP7_75t_R register___U85 ( .A(register__n10785), .Y(register__n5471) );
  CKINVDCx11_ASAP7_75t_R register___U86 ( .A(register__C6422_net59538), .Y(register__n420) );
  AND2x2_ASAP7_75t_R register___U87 ( .A(register__n1514), .B(register__n1515), .Y(register__n20) );
  INVxp67_ASAP7_75t_R register___U88 ( .A(register__n835), .Y(register__n_cell_124812_net160762) );
  INVxp67_ASAP7_75t_R register___U89 ( .A(register__n260), .Y(register__n839) );
  BUFx3_ASAP7_75t_R register___U90 ( .A(register__n3144), .Y(register__n5051) );
  INVx1_ASAP7_75t_R register___U91 ( .A(register__n260), .Y(register__n834) );
  INVx1_ASAP7_75t_R register___U92 ( .A(register__n260), .Y(register__n838) );
  INVx1_ASAP7_75t_R register___U93 ( .A(register__n260), .Y(register__n835) );
  INVx2_ASAP7_75t_R register___U94 ( .A(register__C6422_net60443), .Y(register__n368) );
  INVxp67_ASAP7_75t_R register___U95 ( .A(register__n367), .Y(register__n366) );
  OR2x2_ASAP7_75t_R register___U96 ( .A(register__n11051), .B(register__n11053), .Y(register__n21) );
  AND2x2_ASAP7_75t_R register___U97 ( .A(register__n1840), .B(register__n1841), .Y(register__n22) );
  BUFx10_ASAP7_75t_R register___U98 ( .A(register__net126625), .Y(register__C6422_net70534) );
  INVx3_ASAP7_75t_R register___U99 ( .A(register__C6422_net70534), .Y(register__n1509) );
  OR2x2_ASAP7_75t_R register___U100 ( .A(register__n1978), .B(register__n2635), .Y(register__n23) );
  INVx4_ASAP7_75t_R register___U101 ( .A(register__n1977), .Y(register__n1978) );
  BUFx3_ASAP7_75t_R register___U102 ( .A(register__n4165), .Y(register__n8639) );
  HB1xp67_ASAP7_75t_R register___U103 ( .A(register__n4104), .Y(register__n4103) );
  BUFx2_ASAP7_75t_R register___U104 ( .A(register__n10725), .Y(register__n4245) );
  OR2x2_ASAP7_75t_R register___U105 ( .A(register__n2372), .B(register__n2396), .Y(register__n24) );
  OR2x2_ASAP7_75t_R register___U106 ( .A(register__net100833), .B(register__n1691), .Y(register__n25) );
  OR2x2_ASAP7_75t_R register___U107 ( .A(register__net109852), .B(register__n1691), .Y(register__n26) );
  OR2x2_ASAP7_75t_R register___U108 ( .A(register__n9198), .B(register__n9197), .Y(register__n27) );
  OR3x1_ASAP7_75t_R register___U109 ( .A(register__n252), .B(register__n253), .C(register__n254), .Y(register__n28) );
  OA22x2_ASAP7_75t_R register___U110 ( .A1(register__n1868), .A2(register__n_cell_125487_net184714), .B1(
        n1869), .B2(register__net109643), .Y(register__n29) );
  BUFx16f_ASAP7_75t_R register___U111 ( .A(register__C6422_net60405), .Y(register__n413) );
  BUFx6f_ASAP7_75t_R register___U112 ( .A(register__C6422_net60405), .Y(register__n375) );
  INVx2_ASAP7_75t_R register___U113 ( .A(register__n4710), .Y(register__n8559) );
  INVx1_ASAP7_75t_R register___U114 ( .A(register__n4819), .Y(register__n8248) );
  BUFx2_ASAP7_75t_R register___U115 ( .A(register__n10897), .Y(register__n3141) );
  OR2x2_ASAP7_75t_R register___U116 ( .A(register__n2330), .B(register__n2351), .Y(register__n30) );
  BUFx6f_ASAP7_75t_R register___U117 ( .A(register__net129747), .Y(register__C6422_net70282) );
  INVx3_ASAP7_75t_R register___U118 ( .A(register__C6422_net59572), .Y(register__net129746) );
  BUFx12f_ASAP7_75t_R register___U119 ( .A(register__C6422_net60422), .Y(register__net129747) );
  OR2x2_ASAP7_75t_R register___U120 ( .A(register__n10671), .B(register__n10672), .Y(register__n31) );
  INVx2_ASAP7_75t_R register___U121 ( .A(register__n3097), .Y(register__n7308) );
  INVx2_ASAP7_75t_R register___U122 ( .A(register__n3133), .Y(register__n6451) );
  OR3x1_ASAP7_75t_R register___U123 ( .A(register__n3147), .B(register__n3146), .C(register__n2953), .Y(register__n32) );
  INVx2_ASAP7_75t_R register___U124 ( .A(register__n5062), .Y(register__n7266) );
  INVx1_ASAP7_75t_R register___U125 ( .A(register__n507), .Y(register__n156) );
  INVx3_ASAP7_75t_R register___U126 ( .A(register__n8010), .Y(register__n8012) );
  INVx1_ASAP7_75t_R register___U127 ( .A(register__n3), .Y(register__n158) );
  AO22x1_ASAP7_75t_R register___U128 ( .A1(register__net90661), .A2(register__n3), .B1(register__net89613), .B2(register__n233), 
        .Y(register__n10731) );
  BUFx12f_ASAP7_75t_R register___U129 ( .A(register__n1226), .Y(register__n77) );
  CKINVDCx10_ASAP7_75t_R register___U130 ( .A(register__n11148), .Y(register__n312) );
  BUFx6f_ASAP7_75t_R register___U131 ( .A(register__n381), .Y(register__n281) );
  INVx4_ASAP7_75t_R register___U132 ( .A(register__n2002), .Y(register__n1977) );
  BUFx3_ASAP7_75t_R register___U133 ( .A(register__n2002), .Y(register__n2081) );
  BUFx4f_ASAP7_75t_R register___U134 ( .A(register__n2002), .Y(register__n2080) );
  AND2x6_ASAP7_75t_R register___U135 ( .A(register__n11151), .B(register__n290), .Y(register__net123880) );
  CKINVDCx10_ASAP7_75t_R register___U136 ( .A(register__net96692), .Y(register__n1345) );
  NAND2xp5_ASAP7_75t_R register___U137 ( .A(register__n8783), .B(register__net88727), .Y(register__n349) );
  AND2x6_ASAP7_75t_R register___U138 ( .A(register__n11151), .B(register__n1012), .Y(register__C6422_net59546) );
  CKINVDCx10_ASAP7_75t_R register___U139 ( .A(register__n799), .Y(register__n800) );
  INVx2_ASAP7_75t_R register___U140 ( .A(register__n1993), .Y(register__n1994) );
  OR3x1_ASAP7_75t_R register___U141 ( .A(register__n1032), .B(register__n1033), .C(register__n1034), .Y(register__n11301) );
  NAND2x1p5_ASAP7_75t_R register___U142 ( .A(register__net88752), .B(register__n1993), .Y(register__n2582) );
  INVx6_ASAP7_75t_R register___U143 ( .A(register__n1995), .Y(register__n1993) );
  INVx1_ASAP7_75t_R register___U144 ( .A(register__net112578), .Y(register__n1580) );
  NOR2x2_ASAP7_75t_R register___U145 ( .A(register__n139), .B(register__n724), .Y(register__n768) );
  BUFx4_ASAP7_75t_R register___U146 ( .A(register__n222), .Y(register__n724) );
  NAND2xp5_ASAP7_75t_R register___U147 ( .A(register__n9202), .B(register__n2767), .Y(register__n1501) );
  AO22x2_ASAP7_75t_R register___U148 ( .A1(register__net90237), .A2(register__net109204), .B1(register__net94789), .B2(
        n59), .Y(register__n11092) );
  AO22x2_ASAP7_75t_R register___U149 ( .A1(register__n6975), .A2(register__net109204), .B1(register__n10473), .B2(register__n59), 
        .Y(register__n11050) );
  AO22x2_ASAP7_75t_R register___U150 ( .A1(register__n10436), .A2(register__net109204), .B1(register__n10475), .B2(register__n59), 
        .Y(register__n11073) );
  CKINVDCx10_ASAP7_75t_R register___U151 ( .A(register__net109204), .Y(register__net99656) );
  AO22x2_ASAP7_75t_R register___U152 ( .A1(register__n9670), .A2(register__net109204), .B1(register__n9917), .B2(register__n59), 
        .Y(register__n10945) );
  AO22x2_ASAP7_75t_R register___U153 ( .A1(register__net90853), .A2(register__net109204), .B1(register__net90169), .B2(
        n59), .Y(register__n11008) );
  AO22x2_ASAP7_75t_R register___U154 ( .A1(register__net109204), .A2(register__n9676), .B1(register__n9419), .B2(register__n34), 
        .Y(register__n10608) );
  INVxp67_ASAP7_75t_R register___U155 ( .A(register__n2323), .Y(register__n2348) );
  NOR2x1p5_ASAP7_75t_R register___U156 ( .A(register__C6423_net60623), .B(register__net130087), .Y(register__n2323) );
  AO22x2_ASAP7_75t_R register___U157 ( .A1(register__n7990), .A2(register__C6422_net60422), .B1(register__n9363), .B2(
        net123857), .Y(register__n10671) );
  AO22x2_ASAP7_75t_R register___U158 ( .A1(register__n9605), .A2(register__n39), .B1(register__n10030), .B2(
        C6422_net60399), .Y(register__n10537) );
  AO22x2_ASAP7_75t_R register___U159 ( .A1(register__n9752), .A2(register__n39), .B1(register__n8116), .B2(
        C6422_net60399), .Y(register__n10769) );
  AO22x2_ASAP7_75t_R register___U160 ( .A1(register__n8514), .A2(register__n39), .B1(register__n6662), .B2(
        C6422_net60399), .Y(register__n11024) );
  AO22x2_ASAP7_75t_R register___U161 ( .A1(register__n9814), .A2(register__n39), .B1(register__n8156), .B2(
        C6422_net60399), .Y(register__n10745) );
  AO22x2_ASAP7_75t_R register___U162 ( .A1(register__n9299), .A2(register__n39), .B1(register__n10199), .B2(
        C6422_net60399), .Y(register__n11111) );
  AO22x2_ASAP7_75t_R register___U163 ( .A1(register__n6944), .A2(register__n39), .B1(register__n10241), .B2(
        C6422_net60399), .Y(register__n10896) );
  AO22x2_ASAP7_75t_R register___U164 ( .A1(register__n8795), .A2(register__n39), .B1(register__n8349), .B2(
        C6422_net60399), .Y(register__n10559) );
  BUFx2_ASAP7_75t_R register___U165 ( .A(register__n10718), .Y(register__n4833) );
  INVx1_ASAP7_75t_R register___U166 ( .A(register__n10849), .Y(register__n33) );
  BUFx12f_ASAP7_75t_R register___U167 ( .A(register__n59), .Y(register__n34) );
  BUFx2_ASAP7_75t_R register___U168 ( .A(register__n10929), .Y(register__n4934) );
  BUFx6f_ASAP7_75t_R register___U169 ( .A(register__net123857), .Y(register__net139537) );
  AO22x2_ASAP7_75t_R register___U170 ( .A1(register__n7988), .A2(register__n413), .B1(register__n8799), .B2(register__net126602), 
        .Y(register__n10918) );
  AO22x2_ASAP7_75t_R register___U171 ( .A1(register__n9873), .A2(register__n413), .B1(register__n10287), .B2(register__net126602), 
        .Y(register__n11023) );
  INVx3_ASAP7_75t_R register___U172 ( .A(register__n8012), .Y(register__n1854) );
  INVx1_ASAP7_75t_R register___U173 ( .A(register__n5461), .Y(register__n9231) );
  BUFx2_ASAP7_75t_R register___U174 ( .A(register__n10680), .Y(register__n5461) );
  CKINVDCx11_ASAP7_75t_R register___U175 ( .A(register__C6422_net59548), .Y(register__n817) );
  NOR2x1_ASAP7_75t_R register___U176 ( .A(register__n817), .B(register__n6983), .Y(register__n721) );
  NAND2xp5_ASAP7_75t_R register___U177 ( .A(register__n561), .B(register__n2395), .Y(register__n2394) );
  AND2x6_ASAP7_75t_R register___U178 ( .A(register__n347), .B(register__n312), .Y(register__net119602) );
  INVx6_ASAP7_75t_R register___U179 ( .A(register__n34), .Y(register__n1455) );
  INVx13_ASAP7_75t_R register___U180 ( .A(register__C6422_net59550), .Y(register__net112580) );
  NOR2xp67_ASAP7_75t_R register___U181 ( .A(register__net112580), .B(register__n6469), .Y(register__n622) );
  NOR2x1_ASAP7_75t_R register___U182 ( .A(register__n11183), .B(register__net112580), .Y(register__n722) );
  INVxp67_ASAP7_75t_R register___U183 ( .A(register__n4242), .Y(register__n5520) );
  INVx1_ASAP7_75t_R register___U184 ( .A(register__n11037), .Y(register__n9202) );
  NOR2xp33_ASAP7_75t_R register___U185 ( .A(register__n2347), .B(register__n2322), .Y(register__n2346) );
  NAND2xp5_ASAP7_75t_R register___U186 ( .A(register__n7728), .B(register__n7019), .Y(register__n262) );
  NAND2xp33_ASAP7_75t_R register___U187 ( .A(register__n728), .B(register__n2369), .Y(read_reg_data_1[6]) );
  BUFx16f_ASAP7_75t_R register___U188 ( .A(register__C6422_net60415), .Y(register__net109204) );
  AO22x2_ASAP7_75t_R register___U189 ( .A1(register__n9678), .A2(register__C6422_net60415), .B1(register__n9925), .B2(
        net88727), .Y(register__n10583) );
  NAND2xp67_ASAP7_75t_R register___U190 ( .A(register__n9758), .B(register__C6422_net60415), .Y(register__n256) );
  NAND2xp5_ASAP7_75t_R register___U191 ( .A(register__n49), .B(register__n1501), .Y(register__n556) );
  BUFx2_ASAP7_75t_R register___U192 ( .A(register__n10586), .Y(register__n4449) );
  NAND2xp67_ASAP7_75t_R register___U193 ( .A(register__n9337), .B(register__C6422_net60415), .Y(register__n348) );
  NOR2xp33_ASAP7_75t_R register___U194 ( .A(register__n2665), .B(register__n1892), .Y(register__n2673) );
  AND2x2_ASAP7_75t_R register___U195 ( .A(register__n7321), .B(register__n35), .Y(register__n1882) );
  INVx1_ASAP7_75t_R register___U196 ( .A(register__n10652), .Y(register__n36) );
  AO22x2_ASAP7_75t_R register___U197 ( .A1(register__net90657), .A2(register__n413), .B1(register__net98512), .B2(
        net126602), .Y(register__n10722) );
  AO22x2_ASAP7_75t_R register___U198 ( .A1(register__n8815), .A2(register__net146144), .B1(register__n7221), .B2(
        net126602), .Y(register__n11044) );
  OAI22xp33_ASAP7_75t_R register___U199 ( .A1(register__n53), .A2(register__n7275), .B1(register__net61369), .B2(register__n12327), .Y(read_reg_data_1[20]) );
  AO22x2_ASAP7_75t_R register___U200 ( .A1(register__n9746), .A2(register__C6422_net60405), .B1(register__n8456), .B2(
        C6422_net60401), .Y(register__n10768) );
  AO22x2_ASAP7_75t_R register___U201 ( .A1(register__n9810), .A2(register__C6422_net60405), .B1(register__n10335), .B2(
        C6422_net60401), .Y(register__n11067) );
  AO22x2_ASAP7_75t_R register___U202 ( .A1(register__n9845), .A2(register__C6422_net60405), .B1(register__n6650), .B2(
        C6422_net60401), .Y(register__n10983) );
  AO22x2_ASAP7_75t_R register___U203 ( .A1(register__n9909), .A2(register__n375), .B1(register__n6931), .B2(register__net126602), 
        .Y(register__n11110) );
  HB1xp67_ASAP7_75t_R register___U204 ( .A(register__n10859), .Y(register__n7884) );
  BUFx6f_ASAP7_75t_R register___U205 ( .A(register__net119602), .Y(register__n40) );
  BUFx16f_ASAP7_75t_R register___U206 ( .A(register__net119602), .Y(register__n39) );
  AND2x6_ASAP7_75t_R register___U207 ( .A(register__n11135), .B(register__n312), .Y(register__n799) );
  AND2x6_ASAP7_75t_R register___U208 ( .A(register__n11142), .B(register__n312), .Y(register__n387) );
  INVx3_ASAP7_75t_R register___U209 ( .A(register__net146144), .Y(register__n_cell_125487_net184714) );
  BUFx2_ASAP7_75t_R register___U210 ( .A(register__n2839), .Y(register__n2838) );
  INVxp33_ASAP7_75t_R register___U211 ( .A(register__n155), .Y(register__n37) );
  BUFx12f_ASAP7_75t_R register___U212 ( .A(register__C6422_net60445), .Y(register__n38) );
  NOR4xp25_ASAP7_75t_R register___U213 ( .A(register__n10879), .B(register__n10880), .C(register__n10881), .D(register__n10882), 
        .Y(register__n10859) );
  OAI22xp33_ASAP7_75t_R register___U214 ( .A1(register__n2650), .A2(register__n388), .B1(register__n1455), .B2(register__n2649), 
        .Y(register__n2674) );
  OAI21xp33_ASAP7_75t_R register___U215 ( .A1(register__n2386), .A2(register__n327), .B(register__n2407), .Y(register__n2406) );
  OAI21xp5_ASAP7_75t_R register___U216 ( .A1(register__n2656), .A2(register__n1577), .B(register__n2679), .Y(register__n2680) );
  AO221x2_ASAP7_75t_R register___U217 ( .A1(register__n1361), .A2(register__net91563), .B1(register__n39), .B2(register__net91033), .C(register__n2379), .Y(register__n2398) );
  AO22x1_ASAP7_75t_R register___U218 ( .A1(register__n9662), .A2(register__net104773), .B1(register__n9991), .B2(register__n1350), 
        .Y(register__n10920) );
  NAND2xp5_ASAP7_75t_R register___U219 ( .A(register__n10679), .B(register__n1881), .Y(register__n2162) );
  AND2x6_ASAP7_75t_R register___U220 ( .A(register__n443), .B(register__n11152), .Y(register__C6422_net60437) );
  BUFx6f_ASAP7_75t_R register___U221 ( .A(register__n1345), .Y(register__n41) );
  BUFx12f_ASAP7_75t_R register___U222 ( .A(register__n413), .Y(register__net146144) );
  OAI22xp5_ASAP7_75t_R register___U223 ( .A1(register__n1859), .A2(register__n_cell_125487_net184714), .B1(
        n1860), .B2(register__net109643), .Y(register__n10828) );
  AND2x6_ASAP7_75t_R register___U224 ( .A(register__n443), .B(register__n312), .Y(register__net121619) );
  NAND2x2_ASAP7_75t_R register___U225 ( .A(register__n13), .B(register__n11149), .Y(register__n507) );
  AOI22xp5_ASAP7_75t_R register___U226 ( .A1(register__n9591), .A2(register__net118635), .B1(register__n10012), .B2(
        C6422_net70534), .Y(register__n42) );
  INVx1_ASAP7_75t_R register___U227 ( .A(register__n603), .Y(register__n559) );
  OR2x2_ASAP7_75t_R register___U228 ( .A(register__n2375), .B(register__n1866), .Y(register__n603) );
  INVx1_ASAP7_75t_R register___U229 ( .A(register__net104772), .Y(register__n1866) );
  AND2x2_ASAP7_75t_R register___U230 ( .A(register__n10633), .B(register__n1315), .Y(register__n43) );
  AND3x1_ASAP7_75t_R register___U231 ( .A(register__n43), .B(register__n6142), .C(register__n10635), .Y(register__n8644) );
  BUFx2_ASAP7_75t_R register___U232 ( .A(register__n10634), .Y(register__n6142) );
  AND4x2_ASAP7_75t_R register___U233 ( .A(register__n7936), .B(register__n7934), .C(register__n7935), .D(register__n2205), .Y(
        n10635) );
  BUFx6f_ASAP7_75t_R register___U234 ( .A(register__C6422_net60422), .Y(register__n1853) );
  BUFx3_ASAP7_75t_R register___U235 ( .A(register__net140727), .Y(register__C6422_net59572) );
  INVx2_ASAP7_75t_R register___U236 ( .A(register__C6422_net60422), .Y(register__net140727) );
  OR2x2_ASAP7_75t_R register___U237 ( .A(register__n3525), .B(register__n10806), .Y(register__n44) );
  OR3x2_ASAP7_75t_R register___U238 ( .A(register__n44), .B(register__n10807), .C(register__n1050), .Y(register__n2282) );
  AND3x1_ASAP7_75t_R register___U239 ( .A(register__n6456), .B(register__n6454), .C(register__n6455), .Y(register__n45) );
  AND2x2_ASAP7_75t_R register___U240 ( .A(register__n3372), .B(register__n45), .Y(register__n6453) );
  AND2x2_ASAP7_75t_R register___U241 ( .A(register__n4957), .B(register__C6422_net60405), .Y(register__n46) );
  AND2x2_ASAP7_75t_R register___U242 ( .A(register__n6322), .B(register__C6422_net60401), .Y(register__n47) );
  OR2x2_ASAP7_75t_R register___U243 ( .A(register__n46), .B(register__n47), .Y(register__n10577) );
  BUFx2_ASAP7_75t_R register___U244 ( .A(register__n9331), .Y(register__n4957) );
  BUFx2_ASAP7_75t_R register___U245 ( .A(register__n9357), .Y(register__n6322) );
  NAND2xp5_ASAP7_75t_R register___U246 ( .A(register__n9186), .B(register__n1014), .Y(register__n2160) );
  NAND2xp5_ASAP7_75t_R register___U247 ( .A(register__n1366), .B(register__n1365), .Y(read_reg_data_1[2]) );
  INVx1_ASAP7_75t_R register___U248 ( .A(register__n48), .Y(register__n49) );
  BUFx2_ASAP7_75t_R register___U249 ( .A(register__net61367), .Y(register__n55) );
  AND2x6_ASAP7_75t_R register___U250 ( .A(register__n11141), .B(register__n437), .Y(register__C6422_net60405) );
  OAI21xp33_ASAP7_75t_R register___U251 ( .A1(register__n2410), .A2(register__n2411), .B(register__n51), .Y(register__n2369) );
  AND2x2_ASAP7_75t_R register___U252 ( .A(register__n1760), .B(register__n11150), .Y(register__n56) );
  AND2x6_ASAP7_75t_R register___U253 ( .A(register__n347), .B(register__n13), .Y(register__n1867) );
  INVx1_ASAP7_75t_R register___U254 ( .A(register__n1345), .Y(register__n1361) );
  INVxp67_ASAP7_75t_R register___U255 ( .A(register__n1345), .Y(register__n1344) );
  INVx1_ASAP7_75t_R register___U256 ( .A(register__n1345), .Y(register__n1346) );
  INVx1_ASAP7_75t_R register___U257 ( .A(register__n1345), .Y(register__n1360) );
  INVx1_ASAP7_75t_R register___U258 ( .A(register__n1345), .Y(register__n1359) );
  INVx1_ASAP7_75t_R register___U259 ( .A(register__n1345), .Y(register__n1348) );
  INVxp67_ASAP7_75t_R register___U260 ( .A(register__n1345), .Y(register__n1355) );
  INVx2_ASAP7_75t_R register___U261 ( .A(register__n41), .Y(register__n1347) );
  OR2x2_ASAP7_75t_R register___U262 ( .A(register__n11066), .B(register__n11068), .Y(register__n57) );
  OR3x1_ASAP7_75t_R register___U263 ( .A(register__n57), .B(register__n3497), .C(register__n1375), .Y(register__n64) );
  BUFx2_ASAP7_75t_R register___U264 ( .A(register__n3498), .Y(register__n3497) );
  INVx1_ASAP7_75t_R register___U265 ( .A(register__n1345), .Y(register__n1358) );
  AND2x6_ASAP7_75t_R register___U266 ( .A(register__n11131), .B(register__n11152), .Y(register__C6422_net59542) );
  CKINVDCx11_ASAP7_75t_R register___U267 ( .A(register__C6422_net59542), .Y(register__net107674) );
  AND2x2_ASAP7_75t_R register___U268 ( .A(register__n7149), .B(register__n7646), .Y(register__n58) );
  AND3x1_ASAP7_75t_R register___U269 ( .A(register__n4249), .B(register__n7647), .C(register__n58), .Y(register__n10884) );
  BUFx16f_ASAP7_75t_R register___U270 ( .A(register__net88727), .Y(register__n59) );
  AND2x6_ASAP7_75t_R register___U271 ( .A(register__n11141), .B(register__n11152), .Y(register__net88727) );
  BUFx3_ASAP7_75t_R register___U272 ( .A(register__n59), .Y(register__net129911) );
  AND2x2_ASAP7_75t_R register___U273 ( .A(register__n6718), .B(register__n6829), .Y(register__n60) );
  AND3x1_ASAP7_75t_R register___U274 ( .A(register__n60), .B(register__n4794), .C(register__n6717), .Y(register__n10756) );
  INVx1_ASAP7_75t_R register___U275 ( .A(register__n4795), .Y(register__n6717) );
  AND2x6_ASAP7_75t_R register___U276 ( .A(register__n448), .B(register__n13), .Y(register__C6422_net60422) );
  BUFx6f_ASAP7_75t_R register___U277 ( .A(IF_ID_rs1[3]), .Y(register__n885) );
  AND2x2_ASAP7_75t_R register___U278 ( .A(register__n4909), .B(register__n5666), .Y(register__n61) );
  AND3x1_ASAP7_75t_R register___U279 ( .A(register__n61), .B(register__n8263), .C(register__n8262), .Y(register__n8261) );
  AND3x1_ASAP7_75t_R register___U280 ( .A(register__n8223), .B(register__n8222), .C(register__n5263), .Y(register__n62) );
  AND2x2_ASAP7_75t_R register___U281 ( .A(register__n8224), .B(register__n62), .Y(register__n8221) );
  BUFx4f_ASAP7_75t_R register___U282 ( .A(register__C6422_net60445), .Y(register__net120789) );
  INVx1_ASAP7_75t_R register___U283 ( .A(register__n10713), .Y(register__n63) );
  NOR2xp67_ASAP7_75t_R register___U284 ( .A(register__n64), .B(register__n65), .Y(register__n827) );
  NAND2xp67_ASAP7_75t_R register___U285 ( .A(register__n4569), .B(register__n380), .Y(register__n65) );
  BUFx16f_ASAP7_75t_R register___U286 ( .A(register__net107674), .Y(register__n66) );
  AND2x2_ASAP7_75t_R register___U287 ( .A(register__n42), .B(register__n1267), .Y(register__n67) );
  AND3x1_ASAP7_75t_R register___U288 ( .A(register__n67), .B(register__n4621), .C(register__n1300), .Y(register__n10588) );
  HB1xp67_ASAP7_75t_R register___U289 ( .A(register__n10799), .Y(register__n5308) );
  OR2x6_ASAP7_75t_R register___U290 ( .A(IF_ID_rs1[3]), .B(IF_ID_rs1[4]), .Y(
        n11148) );
  INVx2_ASAP7_75t_R register___U291 ( .A(register__n102), .Y(register__n340) );
  INVx3_ASAP7_75t_R register___U292 ( .A(register__n102), .Y(register__n341) );
  INVx3_ASAP7_75t_R register___U293 ( .A(register__n102), .Y(register__n336) );
  BUFx6f_ASAP7_75t_R register___U294 ( .A(IF_ID_rs1[4]), .Y(register__n11846) );
  BUFx6f_ASAP7_75t_R register___U295 ( .A(register__n11151), .Y(register__n818) );
  AND2x6_ASAP7_75t_R register___U296 ( .A(register__n11151), .B(register__n1760), .Y(register__C6422_net60443) );
  AND2x6_ASAP7_75t_R register___U297 ( .A(IF_ID_rs1[4]), .B(IF_ID_rs1[3]), 
        .Y(register__n11151) );
  AND2x6_ASAP7_75t_R register___U298 ( .A(register__n11135), .B(register__n11151), .Y(register__C6422_net59538) );
  INVx2_ASAP7_75t_R register___U299 ( .A(register__n5721), .Y(register__n11767) );
  INVx4_ASAP7_75t_R register___U300 ( .A(register__n5721), .Y(register__n1415) );
  INVx4_ASAP7_75t_R register___U301 ( .A(register__n5721), .Y(register__n1413) );
  CKINVDCx8_ASAP7_75t_R register___U302 ( .A(register__n102), .Y(register__n337) );
  BUFx12f_ASAP7_75t_R register___U303 ( .A(register__n102), .Y(register__n68) );
  CKINVDCx8_ASAP7_75t_R register___U304 ( .A(register__n12501), .Y(register__n102) );
  INVx6_ASAP7_75t_R register___U305 ( .A(register__n102), .Y(register__n339) );
  AO21x2_ASAP7_75t_R register___U306 ( .A1(register__n326), .A2(register__net89813), .B(register__n2337), .Y(register__n2358) );
  INVx2_ASAP7_75t_R register___U307 ( .A(register__n2358), .Y(register__n69) );
  INVx2_ASAP7_75t_R register___U308 ( .A(register__net61369), .Y(register__n1851) );
  INVx2_ASAP7_75t_R register___U309 ( .A(register__n11301), .Y(register__n70) );
  INVx4_ASAP7_75t_R register___U310 ( .A(register__n3944), .Y(register__n954) );
  INVx4_ASAP7_75t_R register___U311 ( .A(register__n3944), .Y(register__n957) );
  INVx5_ASAP7_75t_R register___U312 ( .A(register__n3944), .Y(register__n953) );
  INVx4_ASAP7_75t_R register___U313 ( .A(register__n3944), .Y(register__n951) );
  INVx5_ASAP7_75t_R register___U314 ( .A(register__n3944), .Y(register__n952) );
  AND2x6_ASAP7_75t_R register___U315 ( .A(register__n1963), .B(register__n796), .Y(register__n3944) );
  AND2x6_ASAP7_75t_R register___U316 ( .A(register__n347), .B(register__n11151), .Y(register__C6422_net60399) );
  BUFx6f_ASAP7_75t_R register___U317 ( .A(register__C6422_net60399), .Y(register__net137523) );
  AND2x6_ASAP7_75t_R register___U318 ( .A(register__n385), .B(register__n830), .Y(register__n12496) );
  CKINVDCx6p67_ASAP7_75t_R register___U319 ( .A(register__n12496), .Y(register__n462) );
  CKINVDCx6p67_ASAP7_75t_R register___U320 ( .A(register__n12496), .Y(register__n459) );
  CKINVDCx6p67_ASAP7_75t_R register___U321 ( .A(register__n12496), .Y(register__n461) );
  OR3x2_ASAP7_75t_R register___U322 ( .A(register__n758), .B(register__n759), .C(register__n760), .Y(register__n11497) );
  INVx2_ASAP7_75t_R register___U323 ( .A(register__n11497), .Y(register__n71) );
  AND2x6_ASAP7_75t_R register___U324 ( .A(register__n10518), .B(register__n12490), .Y(register__n4641) );
  CKINVDCx6p67_ASAP7_75t_R register___U325 ( .A(register__n4641), .Y(register__n578) );
  CKINVDCx6p67_ASAP7_75t_R register___U326 ( .A(register__n4641), .Y(register__n577) );
  CKINVDCx6p67_ASAP7_75t_R register___U327 ( .A(register__n4641), .Y(register__n576) );
  INVx4_ASAP7_75t_R register___U328 ( .A(register__net62822), .Y(register__n72) );
  INVx6_ASAP7_75t_R register___U329 ( .A(register__net124977), .Y(register__net62822) );
  BUFx2_ASAP7_75t_R register___U330 ( .A(register__n7050), .Y(register__n11840) );
  BUFx16f_ASAP7_75t_R register___U331 ( .A(register__n7050), .Y(register__n11843) );
  BUFx3_ASAP7_75t_R register___U332 ( .A(register__n7050), .Y(register__n11838) );
  BUFx16f_ASAP7_75t_R register___U333 ( .A(register__n3280), .Y(register__n12329) );
  BUFx2_ASAP7_75t_R register___U334 ( .A(register__n3280), .Y(register__n12326) );
  BUFx12f_ASAP7_75t_R register___U335 ( .A(register__n3280), .Y(register__n3701) );
  BUFx12f_ASAP7_75t_R register___U336 ( .A(register__n3280), .Y(register__n3702) );
  BUFx16f_ASAP7_75t_R register___U337 ( .A(register__n12336), .Y(register__n3280) );
  NOR2x1p5_ASAP7_75t_R register___U338 ( .A(register__n9363), .B(register__n1473), .Y(register__n2792) );
  BUFx4f_ASAP7_75t_R register___U339 ( .A(register__n3021), .Y(register__n1473) );
  BUFx10_ASAP7_75t_R register___U340 ( .A(register__n12498), .Y(register__n1887) );
  OR2x2_ASAP7_75t_R register___U341 ( .A(register__n8710), .B(register__n2818), .Y(register__n2796) );
  INVx3_ASAP7_75t_R register___U342 ( .A(register__n2796), .Y(register__n73) );
  NOR2xp67_ASAP7_75t_R register___U343 ( .A(register__C6423_net72545), .B(register__n1886), .Y(register__n2525) );
  AND2x4_ASAP7_75t_R register___U344 ( .A(register__n11714), .B(register__n7052), .Y(register__n11729) );
  BUFx2_ASAP7_75t_R register___U345 ( .A(rs2[1]), .Y(register__n2233) );
  BUFx4f_ASAP7_75t_R register___U346 ( .A(rs2[1]), .Y(register__n406) );
  NOR2x1p5_ASAP7_75t_R register___U347 ( .A(register__n11726), .B(register__n2739), .Y(register__net93897) );
  BUFx12f_ASAP7_75t_R register___U348 ( .A(register__net130482), .Y(register__net141879) );
  HB1xp67_ASAP7_75t_R register___U349 ( .A(register__net130482), .Y(register__net66614) );
  BUFx4f_ASAP7_75t_R register___U350 ( .A(register__net130482), .Y(register__net66618) );
  OAI22xp5_ASAP7_75t_R register___U351 ( .A1(register__net66314), .A2(register__n8272), .B1(register__n5345), .B2(register__n1687), .Y(read_reg_data_2[21]) );
  AND3x1_ASAP7_75t_R register___U352 ( .A(register__n843), .B(register__n9241), .C(register__n11542), .Y(register__n8272) );
  INVx1_ASAP7_75t_R register___U353 ( .A(register__n11544), .Y(register__n5994) );
  INVx4_ASAP7_75t_R register___U354 ( .A(rs2[0]), .Y(register__n11721) );
  INVx2_ASAP7_75t_R register___U355 ( .A(register__n11709), .Y(register__n2222) );
  INVx1_ASAP7_75t_R register___U356 ( .A(register__n264), .Y(register__n601) );
  INVx1_ASAP7_75t_R register___U357 ( .A(register__n5441), .Y(register__n264) );
  BUFx4f_ASAP7_75t_R register___U358 ( .A(rs2[0]), .Y(register__n2277) );
  AOI211xp5_ASAP7_75t_R register___U359 ( .A1(register__n650), .A2(register__net89397), .B(register__n2735), .C(register__n2737), 
        .Y(register__n2738) );
  BUFx6f_ASAP7_75t_R register___U360 ( .A(rs2[2]), .Y(register__n5441) );
  INVx4_ASAP7_75t_R register___U361 ( .A(register__n1129), .Y(register__n_cell_125074_net170554) );
  NOR3xp33_ASAP7_75t_R register___U362 ( .A(register__n287), .B(register__n1167), .C(register__n1166), .Y(register__n11540) );
  INVxp67_ASAP7_75t_R register___U363 ( .A(register__n286), .Y(register__n287) );
  AO22x2_ASAP7_75t_R register___U364 ( .A1(register__n10509), .A2(register__net110414), .B1(register__n10511), .B2(
        net125797), .Y(register__n11557) );
  NOR2x2_ASAP7_75t_R register___U365 ( .A(register__n1036), .B(register__n11727), .Y(register__n1129) );
  NOR2x1p5_ASAP7_75t_R register___U366 ( .A(register__n8783), .B(register__n1629), .Y(register__n2783) );
  INVx3_ASAP7_75t_R register___U367 ( .A(register__n3268), .Y(register__n1629) );
  INVx1_ASAP7_75t_R register___U368 ( .A(register__n5460), .Y(register__n1041) );
  INVx1_ASAP7_75t_R register___U369 ( .A(register__net130482), .Y(register__n2118) );
  INVx2_ASAP7_75t_R register___U370 ( .A(register__net130482), .Y(register__n2119) );
  INVx2_ASAP7_75t_R register___U371 ( .A(register__net130482), .Y(register__n2117) );
  INVx2_ASAP7_75t_R register___U372 ( .A(register__net130482), .Y(register__n1653) );
  CKINVDCx10_ASAP7_75t_R register___U373 ( .A(register__n488), .Y(register__n422) );
  AND4x2_ASAP7_75t_R register___U374 ( .A(register__n9173), .B(register__n3699), .C(register__n9172), .D(register__n2997), .Y(
        n159) );
  INVx2_ASAP7_75t_R register___U375 ( .A(register__n159), .Y(register__n74) );
  INVx2_ASAP7_75t_R register___U376 ( .A(register__n5212), .Y(register__n1557) );
  INVx1_ASAP7_75t_R register___U377 ( .A(register__n2883), .Y(register__n1806) );
  INVx1_ASAP7_75t_R register___U378 ( .A(register__n4756), .Y(register__n1068) );
  INVx3_ASAP7_75t_R register___U379 ( .A(register__net112585), .Y(register__C6422_net59961) );
  BUFx16f_ASAP7_75t_R register___U380 ( .A(register__C6422_net60437), .Y(register__n75) );
  AND2x4_ASAP7_75t_R register___U381 ( .A(register__net125365), .B(register__net89010), .Y(register__n2570) );
  INVx2_ASAP7_75t_R register___U382 ( .A(register__n2570), .Y(register__n76) );
  INVx1_ASAP7_75t_R register___U383 ( .A(register__n11204), .Y(register__n247) );
  NAND2x2_ASAP7_75t_R register___U384 ( .A(register__n334), .B(register__net89661), .Y(register__n2627) );
  AND2x6_ASAP7_75t_R register___U385 ( .A(register__n11720), .B(register__n11728), .Y(register__n334) );
  INVx2_ASAP7_75t_R register___U386 ( .A(register__n9636), .Y(register__n1759) );
  INVx1_ASAP7_75t_R register___U387 ( .A(register__n9636), .Y(register__n1859) );
  AO22x2_ASAP7_75t_R register___U388 ( .A1(register__n9636), .A2(register__net125170), .B1(register__n9421), .B2(register__n515), 
        .Y(register__n11438) );
  INVx2_ASAP7_75t_R register___U389 ( .A(register__n9949), .Y(register__n664) );
  INVx3_ASAP7_75t_R register___U390 ( .A(register__C6423_net61318), .Y(register__net126725) );
  INVx2_ASAP7_75t_R register___U391 ( .A(register__C6423_net61318), .Y(register__n1172) );
  INVx2_ASAP7_75t_R register___U392 ( .A(register__C6423_net61318), .Y(register__n1171) );
  AO22x1_ASAP7_75t_R register___U393 ( .A1(register__net63216), .A2(register__n342), .B1(register__n1877), .B2(register__n339), 
        .Y(register__n1876) );
  AO22x1_ASAP7_75t_R register___U394 ( .A1(register__net139893), .A2(register__n1590), .B1(register__net105510), .B2(
        n3022), .Y(register__n736) );
  AO22x1_ASAP7_75t_R register___U395 ( .A1(register__net140270), .A2(register__n1058), .B1(register__net105518), .B2(
        n1140), .Y(register__n1008) );
  AO22x1_ASAP7_75t_R register___U396 ( .A1(register__net63362), .A2(register__n1306), .B1(register__n1307), .B2(register__n1308), 
        .Y(register__n1305) );
  NOR4xp25_ASAP7_75t_R register___U397 ( .A(register__n2535), .B(register__n2534), .C(register__n2533), .D(register__n2561), .Y(
        n2560) );
  NOR2xp67_ASAP7_75t_R register___U398 ( .A(register__net105488), .B(register__n711), .Y(register__n2535) );
  AO22x1_ASAP7_75t_R register___U399 ( .A1(register__net64868), .A2(register__n896), .B1(register__n1426), .B2(register__n889), 
        .Y(register__n1425) );
  BUFx2_ASAP7_75t_R register___U400 ( .A(register__n12250), .Y(register__n733) );
  BUFx8_ASAP7_75t_R register___U401 ( .A(register__n12250), .Y(register__n12249) );
  BUFx2_ASAP7_75t_R register___U402 ( .A(register__n12250), .Y(register__n732) );
  INVx2_ASAP7_75t_R register___U403 ( .A(register__n4968), .Y(register__n1861) );
  INVx4_ASAP7_75t_R register___U404 ( .A(register__n4968), .Y(register__n889) );
  INVx4_ASAP7_75t_R register___U405 ( .A(register__n4968), .Y(register__n895) );
  INVx4_ASAP7_75t_R register___U406 ( .A(register__n4968), .Y(register__n894) );
  INVx4_ASAP7_75t_R register___U407 ( .A(register__n4968), .Y(register__n893) );
  INVx5_ASAP7_75t_R register___U408 ( .A(register__n4968), .Y(register__n890) );
  AND2x6_ASAP7_75t_R register___U409 ( .A(register__n1963), .B(register__n3407), .Y(register__n4968) );
  OA21x2_ASAP7_75t_R register___U410 ( .A1(register__net105496), .A2(register__n712), .B(register__n2444), .Y(register__n2445) );
  INVx3_ASAP7_75t_R register___U411 ( .A(register__n2445), .Y(register__n78) );
  NOR2x1p5_ASAP7_75t_R register___U412 ( .A(register__n406), .B(register__n79), .Y(register__n1107) );
  NOR2x2_ASAP7_75t_R register___U413 ( .A(register__n430), .B(register__n5441), .Y(register__n80) );
  INVx2_ASAP7_75t_R register___U414 ( .A(register__n80), .Y(register__n79) );
  BUFx6f_ASAP7_75t_R register___U415 ( .A(rs2[0]), .Y(register__n430) );
  BUFx24_ASAP7_75t_R register___U416 ( .A(register__n5720), .Y(register__n81) );
  BUFx24_ASAP7_75t_R register___U417 ( .A(register__n5720), .Y(register__n82) );
  INVxp67_ASAP7_75t_R register___U418 ( .A(register__n1313), .Y(register__n1493) );
  NOR2xp67_ASAP7_75t_R register___U419 ( .A(register__n1314), .B(register__n_cell_125074_net170554), .Y(register__n1313) );
  INVx1_ASAP7_75t_R register___U420 ( .A(register__n1887), .Y(register__n2827) );
  INVx1_ASAP7_75t_R register___U421 ( .A(register__n1887), .Y(register__n2824) );
  INVx1_ASAP7_75t_R register___U422 ( .A(register__n1887), .Y(register__n2822) );
  INVx1_ASAP7_75t_R register___U423 ( .A(register__n1887), .Y(register__n2823) );
  INVx1_ASAP7_75t_R register___U424 ( .A(register__n1887), .Y(register__n2825) );
  INVx6_ASAP7_75t_R register___U425 ( .A(register__n1652), .Y(register__n111) );
  BUFx12f_ASAP7_75t_R register___U426 ( .A(register__net130482), .Y(register__n1652) );
  CKINVDCx6p67_ASAP7_75t_R register___U427 ( .A(register__n1656), .Y(register__n110) );
  BUFx12f_ASAP7_75t_R register___U428 ( .A(register__net130482), .Y(register__n1656) );
  INVx6_ASAP7_75t_R register___U429 ( .A(register__net123862), .Y(register__n112) );
  BUFx12f_ASAP7_75t_R register___U430 ( .A(register__C6423_net61340), .Y(register__net123862) );
  BUFx3_ASAP7_75t_R register___U431 ( .A(register__n11154), .Y(register__n139) );
  BUFx12f_ASAP7_75t_R register___U432 ( .A(register__n12249), .Y(register__n12245) );
  NAND2xp5_ASAP7_75t_R register___U433 ( .A(register__n6605), .B(register__net88572), .Y(register__n862) );
  BUFx16f_ASAP7_75t_R register___U434 ( .A(register__C6422_net60408), .Y(register__net117658) );
  NOR2x1p5_ASAP7_75t_R register___U435 ( .A(register__n1036), .B(register__n11727), .Y(register__n1073) );
  OR3x4_ASAP7_75t_R register___U436 ( .A(register__n2222), .B(register__n601), .C(register__n2277), .Y(register__n11727) );
  CKINVDCx6p67_ASAP7_75t_R register___U437 ( .A(register__n2141), .Y(register__n1922) );
  INVx5_ASAP7_75t_R register___U438 ( .A(register__n118), .Y(register__n2141) );
  CKINVDCx5p33_ASAP7_75t_R register___U439 ( .A(register__n1049), .Y(register__n3338) );
  CKINVDCx12_ASAP7_75t_R register___U440 ( .A(register__n3276), .Y(register__n1049) );
  OAI22x1_ASAP7_75t_R register___U441 ( .A1(register__net64668), .A2(register__n1049), .B1(register__n6631), .B2(register__n2881), 
        .Y(register__n501) );
  AO22x2_ASAP7_75t_R register___U442 ( .A1(register__net140270), .A2(register__n11751), .B1(register__n2594), .B2(register__n1049), .Y(register__n825) );
  INVx6_ASAP7_75t_R register___U443 ( .A(register__n5721), .Y(register__n1416) );
  AND2x6_ASAP7_75t_R register___U444 ( .A(register__n12492), .B(register__n12490), .Y(register__n5721) );
  INVx1_ASAP7_75t_R register___U445 ( .A(register__n4035), .Y(register__n1591) );
  BUFx4f_ASAP7_75t_R register___U446 ( .A(register__n4035), .Y(register__n4269) );
  INVx6_ASAP7_75t_R register___U447 ( .A(register__n3190), .Y(register__n4035) );
  CKINVDCx20_ASAP7_75t_R register___U448 ( .A(register__n1164), .Y(register__n11730) );
  BUFx24_ASAP7_75t_R register___U449 ( .A(register__n4127), .Y(register__n1164) );
  CKINVDCx10_ASAP7_75t_R register___U450 ( .A(register__n1655), .Y(register__n117) );
  BUFx16f_ASAP7_75t_R register___U451 ( .A(register__net130482), .Y(register__n1655) );
  BUFx12f_ASAP7_75t_R register___U452 ( .A(register__net130482), .Y(register__n1654) );
  AND2x6_ASAP7_75t_R register___U453 ( .A(register__n12484), .B(register__n1904), .Y(register__net130482) );
  INVx5_ASAP7_75t_R register___U454 ( .A(register__n5548), .Y(register__n1647) );
  INVx1_ASAP7_75t_R register___U455 ( .A(register__n1793), .Y(register__n1622) );
  OAI22x1_ASAP7_75t_R register___U456 ( .A1(register__n12152), .A2(register__n1647), .B1(register__n6113), .B2(register__n1640), 
        .Y(register__n706) );
  INVx4_ASAP7_75t_R register___U457 ( .A(register__n5548), .Y(register__n1793) );
  INVx2_ASAP7_75t_R register___U458 ( .A(register__n1792), .Y(register__n1620) );
  NOR2x2_ASAP7_75t_R register___U459 ( .A(register__n9951), .B(register__n82), .Y(register__n8600) );
  AOI22x1_ASAP7_75t_R register___U460 ( .A1(register__net64390), .A2(register__n82), .B1(register__n227), .B2(register__n665), 
        .Y(register__n12820) );
  CKINVDCx11_ASAP7_75t_R register___U461 ( .A(register__net109611), .Y(register__n1987) );
  BUFx2_ASAP7_75t_R register___U462 ( .A(register__n4166), .Y(register__n4165) );
  INVx4_ASAP7_75t_R register___U463 ( .A(register__net93897), .Y(register__n83) );
  INVx3_ASAP7_75t_R register___U464 ( .A(register__n83), .Y(register__n84) );
  INVx5_ASAP7_75t_R register___U465 ( .A(register__n83), .Y(register__n85) );
  BUFx6f_ASAP7_75t_R register___U466 ( .A(register__n11759), .Y(register__n3675) );
  BUFx12f_ASAP7_75t_R register___U467 ( .A(register__n3476), .Y(register__n6430) );
  INVxp67_ASAP7_75t_R register___U468 ( .A(register__n1816), .Y(register__n990) );
  INVxp67_ASAP7_75t_R register___U469 ( .A(register__n5516), .Y(register__n989) );
  BUFx4_ASAP7_75t_R register___U470 ( .A(register__n4636), .Y(register__n12127) );
  INVx3_ASAP7_75t_R register___U471 ( .A(register__n4633), .Y(register__n12120) );
  BUFx10_ASAP7_75t_R register___U472 ( .A(register__n4636), .Y(register__n12128) );
  INVx2_ASAP7_75t_R register___U473 ( .A(register__n12128), .Y(register__n12111) );
  OR2x4_ASAP7_75t_R register___U474 ( .A(register__n1335), .B(register__n7697), .Y(register__n276) );
  INVx1_ASAP7_75t_R register___U475 ( .A(register__n11345), .Y(register__n773) );
  AND2x6_ASAP7_75t_R register___U476 ( .A(register__n7020), .B(register__n11729), .Y(register__C6423_net61318) );
  AND2x6_ASAP7_75t_R register___U477 ( .A(register__n11728), .B(register__n11729), .Y(register__net94400) );
  AND2x6_ASAP7_75t_R register___U478 ( .A(register__n877), .B(register__n11728), .Y(register__C6423_net61348) );
  CKINVDCx5p33_ASAP7_75t_R register___U479 ( .A(register__n651), .Y(register__C6423_net61343) );
  BUFx3_ASAP7_75t_R register___U480 ( .A(register__C6423_net61343), .Y(register__net104685) );
  AO22x1_ASAP7_75t_R register___U481 ( .A1(register__n9575), .A2(register__C6423_net61326), .B1(register__n9431), .B2(
        n2001), .Y(register__n11207) );
  BUFx4f_ASAP7_75t_R register___U482 ( .A(register__C6423_net61326), .Y(register__C6423_net68950) );
  AND2x6_ASAP7_75t_R register___U483 ( .A(register__n11719), .B(register__n11728), .Y(register__n767) );
  AND2x6_ASAP7_75t_R register___U484 ( .A(rs2[3]), .B(register__n8835), .Y(register__n11728) );
  INVx2_ASAP7_75t_R register___U485 ( .A(rs2[4]), .Y(register__n8835) );
  OR3x2_ASAP7_75t_R register___U486 ( .A(register__n428), .B(register__n11143), .C(IF_ID_rs1[2]), .Y(
        n11154) );
  AND2x6_ASAP7_75t_R register___U487 ( .A(register__n347), .B(register__n13), .Y(register__net91683) );
  AND2x6_ASAP7_75t_R register___U488 ( .A(register__n11131), .B(register__n437), .Y(register__C6422_net59550) );
  AND2x4_ASAP7_75t_R register___U489 ( .A(register__n4490), .B(register__n11136), .Y(register__n347) );
  BUFx2_ASAP7_75t_R register___U490 ( .A(register__n10802), .Y(register__n5157) );
  BUFx4f_ASAP7_75t_R register___U491 ( .A(IF_ID_rs1[0]), .Y(register__n11143) );
  NOR2xp33_ASAP7_75t_R register___U492 ( .A(register__n2749), .B(register__n2748), .Y(register__n86) );
  NOR2xp33_ASAP7_75t_R register___U493 ( .A(register__n2747), .B(register__n87), .Y(register__n6019) );
  INVxp33_ASAP7_75t_R register___U494 ( .A(register__n86), .Y(register__n87) );
  NOR2xp33_ASAP7_75t_R register___U495 ( .A(register__n1995), .B(register__net113157), .Y(register__n2748) );
  NOR2xp33_ASAP7_75t_R register___U496 ( .A(register__n1800), .B(register__n5245), .Y(register__n2749) );
  BUFx12f_ASAP7_75t_R register___U497 ( .A(register__n608), .Y(register__n12075) );
  INVx4_ASAP7_75t_R register___U498 ( .A(n4), .Y(register__n608) );
  BUFx4_ASAP7_75t_R register___U499 ( .A(register__n608), .Y(register__n12065) );
  INVx3_ASAP7_75t_R register___U500 ( .A(register__n608), .Y(register__n12051) );
  BUFx10_ASAP7_75t_R register___U501 ( .A(register__n608), .Y(register__n12066) );
  INVxp67_ASAP7_75t_R register___U502 ( .A(register__n2907), .Y(register__n3873) );
  BUFx5_ASAP7_75t_R register___U503 ( .A(register__n12499), .Y(register__n3021) );
  BUFx6f_ASAP7_75t_R register___U504 ( .A(register__n3908), .Y(register__n3909) );
  BUFx16f_ASAP7_75t_R register___U505 ( .A(register__n3908), .Y(register__n11752) );
  INVxp67_ASAP7_75t_R register___U506 ( .A(register__n1836), .Y(register__n88) );
  INVx2_ASAP7_75t_R register___U507 ( .A(register__n1836), .Y(register__n1696) );
  INVx2_ASAP7_75t_R register___U508 ( .A(register__n1836), .Y(register__n1695) );
  INVx2_ASAP7_75t_R register___U509 ( .A(register__n1836), .Y(register__n1692) );
  BUFx3_ASAP7_75t_R register___U510 ( .A(register__n1695), .Y(register__n4575) );
  BUFx4_ASAP7_75t_R register___U511 ( .A(register__n1694), .Y(register__n6160) );
  BUFx8_ASAP7_75t_R register___U512 ( .A(register__n1695), .Y(register__n3354) );
  INVx1_ASAP7_75t_R register___U513 ( .A(register__n1716), .Y(register__n1717) );
  BUFx3_ASAP7_75t_R register___U514 ( .A(register__n1112), .Y(register__n5170) );
  BUFx12f_ASAP7_75t_R register___U515 ( .A(register__n3354), .Y(register__n3353) );
  BUFx4f_ASAP7_75t_R register___U516 ( .A(register__n11871), .Y(register__n3418) );
  INVx1_ASAP7_75t_R register___U517 ( .A(register__n1738), .Y(register__n1739) );
  BUFx6f_ASAP7_75t_R register___U518 ( .A(register__n11871), .Y(register__n11753) );
  BUFx2_ASAP7_75t_R register___U519 ( .A(register__n5170), .Y(register__n11870) );
  INVxp67_ASAP7_75t_R register___U520 ( .A(register__n1730), .Y(register__n1731) );
  BUFx6f_ASAP7_75t_R register___U521 ( .A(register__n11753), .Y(register__n3681) );
  BUFx2_ASAP7_75t_R register___U522 ( .A(register__n11870), .Y(register__n11872) );
  BUFx2_ASAP7_75t_R register___U523 ( .A(register__n11870), .Y(register__n3419) );
  INVxp33_ASAP7_75t_R register___U524 ( .A(register__n1733), .Y(register__n1734) );
  OR2x4_ASAP7_75t_R register___U525 ( .A(register__n2167), .B(register__n1503), .Y(register__n1836) );
  INVx1_ASAP7_75t_R register___U526 ( .A(register__n1696), .Y(register__n1713) );
  INVx1_ASAP7_75t_R register___U527 ( .A(register__n1695), .Y(register__n1705) );
  INVx1_ASAP7_75t_R register___U528 ( .A(register__n1692), .Y(register__n1704) );
  INVx1_ASAP7_75t_R register___U529 ( .A(register__n1692), .Y(register__n1701) );
  INVxp67_ASAP7_75t_R register___U530 ( .A(register__n1696), .Y(register__n1698) );
  INVx1_ASAP7_75t_R register___U531 ( .A(register__n1692), .Y(register__n1716) );
  INVx2_ASAP7_75t_R register___U532 ( .A(register__n1694), .Y(register__n1707) );
  INVx1_ASAP7_75t_R register___U533 ( .A(register__n1692), .Y(register__n1711) );
  INVx2_ASAP7_75t_R register___U534 ( .A(register__n1695), .Y(register__n1720) );
  INVxp67_ASAP7_75t_R register___U535 ( .A(register__n1696), .Y(register__n1712) );
  INVx1_ASAP7_75t_R register___U536 ( .A(register__n1696), .Y(register__n1702) );
  INVx1_ASAP7_75t_R register___U537 ( .A(register__n1695), .Y(register__n1699) );
  INVx1_ASAP7_75t_R register___U538 ( .A(register__n1695), .Y(register__n1703) );
  INVx1_ASAP7_75t_R register___U539 ( .A(register__n1696), .Y(register__n1710) );
  INVx1_ASAP7_75t_R register___U540 ( .A(register__n1692), .Y(register__n1714) );
  INVx1_ASAP7_75t_R register___U541 ( .A(register__n1696), .Y(register__n1706) );
  INVx1_ASAP7_75t_R register___U542 ( .A(register__n1692), .Y(register__n1700) );
  INVxp67_ASAP7_75t_R register___U543 ( .A(register__n1697), .Y(register__n1709) );
  INVx1_ASAP7_75t_R register___U544 ( .A(register__n6160), .Y(register__n1724) );
  INVx1_ASAP7_75t_R register___U545 ( .A(register__n1721), .Y(register__n1722) );
  INVx2_ASAP7_75t_R register___U546 ( .A(register__n4575), .Y(register__n1718) );
  INVx2_ASAP7_75t_R register___U547 ( .A(register__n11871), .Y(register__n1725) );
  INVx3_ASAP7_75t_R register___U548 ( .A(register__n3352), .Y(register__n1736) );
  INVx1_ASAP7_75t_R register___U549 ( .A(register__n1715), .Y(register__n1735) );
  INVx2_ASAP7_75t_R register___U550 ( .A(register__n5170), .Y(register__n1730) );
  INVx1_ASAP7_75t_R register___U551 ( .A(register__n11753), .Y(register__n1729) );
  INVx2_ASAP7_75t_R register___U552 ( .A(register__n3418), .Y(register__n1727) );
  INVx2_ASAP7_75t_R register___U553 ( .A(register__n11870), .Y(register__n1733) );
  INVx2_ASAP7_75t_R register___U554 ( .A(register__n3681), .Y(register__n1732) );
  INVxp67_ASAP7_75t_R register___U555 ( .A(register__n5765), .Y(register__n7033) );
  OR2x4_ASAP7_75t_R register___U556 ( .A(register__n12491), .B(register__n2127), .Y(register__n12501) );
  NAND2xp5_ASAP7_75t_R register___U557 ( .A(register__n51), .B(register__n605), .Y(register__n242) );
  NAND2xp5_ASAP7_75t_R register___U558 ( .A(register__n12), .B(register__n360), .Y(register__n605) );
  INVx3_ASAP7_75t_R register___U559 ( .A(register__n1092), .Y(register__n417) );
  NAND2xp5_ASAP7_75t_R register___U560 ( .A(register__n12485), .B(register__n12503), .Y(register__n594) );
  BUFx2_ASAP7_75t_R register___U561 ( .A(register__n12505), .Y(register__n7678) );
  BUFx6f_ASAP7_75t_R register___U562 ( .A(WB_rd[0]), .Y(register__n1128) );
  BUFx6f_ASAP7_75t_R register___U563 ( .A(register__net147907), .Y(register__net148003) );
  INVx13_ASAP7_75t_R register___U564 ( .A(register__n1975), .Y(register__n1972) );
  BUFx12f_ASAP7_75t_R register___U565 ( .A(register__n2843), .Y(register__n2135) );
  BUFx6f_ASAP7_75t_R register___U566 ( .A(WB_rd[2]), .Y(register__n154) );
  INVx2_ASAP7_75t_R register___U567 ( .A(register__n3408), .Y(register__n1131) );
  INVx3_ASAP7_75t_R register___U568 ( .A(register__n1836), .Y(register__n1694) );
  BUFx12f_ASAP7_75t_R register___U569 ( .A(register__net64038), .Y(register__net64052) );
  BUFx12f_ASAP7_75t_R register___U570 ( .A(register__net142400), .Y(register__net64038) );
  AOI22x1_ASAP7_75t_R register___U571 ( .A1(register__n3531), .A2(register__net130482), .B1(register__n663), .B2(
        net66574), .Y(register__n12638) );
  BUFx6f_ASAP7_75t_R register___U572 ( .A(register__n6139), .Y(register__n4842) );
  BUFx3_ASAP7_75t_R register___U573 ( .A(register__n1510), .Y(register__n4841) );
  CKINVDCx10_ASAP7_75t_R register___U574 ( .A(register__n12125), .Y(register__n6680) );
  BUFx4f_ASAP7_75t_R register___U575 ( .A(register__n12132), .Y(register__n12136) );
  INVx1_ASAP7_75t_R register___U576 ( .A(register__n12136), .Y(register__n12117) );
  BUFx4_ASAP7_75t_R register___U577 ( .A(register__n12497), .Y(register__n2843) );
  CKINVDCx12_ASAP7_75t_R register___U578 ( .A(register__n1972), .Y(register__n1973) );
  BUFx3_ASAP7_75t_R register___U579 ( .A(register__n11798), .Y(register__n11795) );
  INVx2_ASAP7_75t_R register___U580 ( .A(register__n7327), .Y(register__n89) );
  INVx11_ASAP7_75t_R register___U581 ( .A(register__n12504), .Y(register__n7327) );
  BUFx3_ASAP7_75t_R register___U582 ( .A(register__n5788), .Y(register__n5787) );
  INVx1_ASAP7_75t_R register___U583 ( .A(register__n1345), .Y(register__n90) );
  INVx1_ASAP7_75t_R register___U584 ( .A(register__n1345), .Y(register__n91) );
  AND2x6_ASAP7_75t_R register___U585 ( .A(register__n11135), .B(register__n11152), .Y(register__net96692) );
  INVx1_ASAP7_75t_R register___U586 ( .A(register__n1345), .Y(register__n1357) );
  INVx1_ASAP7_75t_R register___U587 ( .A(register__n1345), .Y(register__n1356) );
  INVx1_ASAP7_75t_R register___U588 ( .A(register__n1345), .Y(register__n1354) );
  INVx1_ASAP7_75t_R register___U589 ( .A(register__n1345), .Y(register__n1352) );
  INVx1_ASAP7_75t_R register___U590 ( .A(register__n1345), .Y(register__n1349) );
  BUFx6f_ASAP7_75t_R register___U591 ( .A(register__net64478), .Y(register__net64476) );
  BUFx16f_ASAP7_75t_R register___U592 ( .A(register__n11732), .Y(register__n11731) );
  BUFx12f_ASAP7_75t_R register___U593 ( .A(register__n5182), .Y(register__n11732) );
  BUFx16f_ASAP7_75t_R register___U594 ( .A(register__n6721), .Y(register__n5182) );
  INVxp67_ASAP7_75t_R register___U595 ( .A(register__n3781), .Y(register__n5241) );
  CKINVDCx10_ASAP7_75t_R register___U596 ( .A(WB_rd[0]), .Y(register__n12488) );
  CKINVDCx5p33_ASAP7_75t_R register___U597 ( .A(write_data[15]), .Y(register__net142400) );
  AND2x6_ASAP7_75t_R register___U598 ( .A(register__n347), .B(register__n11152), .Y(register__C6422_net60401) );
  AND2x6_ASAP7_75t_R register___U599 ( .A(register__n726), .B(register__n11152), .Y(register__n381) );
  BUFx3_ASAP7_75t_R register___U600 ( .A(register__n2940), .Y(register__n2939) );
  CKINVDCx16_ASAP7_75t_R register___U601 ( .A(register__n2891), .Y(register__n1975) );
  BUFx2_ASAP7_75t_R register___U602 ( .A(register__n6266), .Y(register__n12436) );
  BUFx12f_ASAP7_75t_R register___U603 ( .A(register__n12504), .Y(register__n5172) );
  OAI22xp5_ASAP7_75t_R register___U604 ( .A1(register__n12236), .A2(register__n7327), .B1(register__n8347), .B2(register__n5172), 
        .Y(register__n408) );
  INVx2_ASAP7_75t_R register___U605 ( .A(register__n5172), .Y(register__n1403) );
  INVx3_ASAP7_75t_R register___U606 ( .A(register__n3572), .Y(register__n1616) );
  INVxp67_ASAP7_75t_R register___U607 ( .A(register__n1160), .Y(register__n775) );
  BUFx8_ASAP7_75t_R register___U608 ( .A(register__net91939), .Y(register__net64452) );
  BUFx4_ASAP7_75t_R register___U609 ( .A(register__n6139), .Y(register__n11904) );
  AOI22xp5_ASAP7_75t_R register___U610 ( .A1(register__n12412), .A2(register__n1972), .B1(register__n523), .B2(register__n524), 
        .Y(register__n12893) );
  CKINVDCx11_ASAP7_75t_R register___U611 ( .A(register__n2135), .Y(register__n1974) );
  AND2x6_ASAP7_75t_R register___U612 ( .A(register__n10518), .B(register__n7684), .Y(register__n6721) );
  INVx2_ASAP7_75t_R register___U613 ( .A(register__n4631), .Y(register__n11876) );
  NAND2xp33_ASAP7_75t_R register___U614 ( .A(register__n1343), .B(register__n2634), .Y(read_reg_data_1[24])
         );
  BUFx6f_ASAP7_75t_R register___U615 ( .A(register__net62718), .Y(register__net62680) );
  INVx4_ASAP7_75t_R register___U616 ( .A(write_data[31]), .Y(register__net62718) );
  NOR2xp67_ASAP7_75t_R register___U617 ( .A(register__n2161), .B(register__n2162), .Y(register__n7939) );
  AOI22xp5_ASAP7_75t_R register___U618 ( .A1(register__net64446), .A2(register__n879), .B1(register__n880), .B2(
        net67384), .Y(register__n13105) );
  BUFx3_ASAP7_75t_R register___U619 ( .A(register__n3328), .Y(register__n11902) );
  BUFx4f_ASAP7_75t_R register___U620 ( .A(register__n12130), .Y(register__n3628) );
  INVx4_ASAP7_75t_R register___U621 ( .A(write_data[12]), .Y(register__n12141) );
  INVx1_ASAP7_75t_R register___U622 ( .A(register__n13026), .Y(register__n92) );
  INVx2_ASAP7_75t_R register___U623 ( .A(register__n12120), .Y(register__n554) );
  BUFx4f_ASAP7_75t_R register___U624 ( .A(register__n1129), .Y(register__net117890) );
  INVx1_ASAP7_75t_R register___U625 ( .A(register__n1707), .Y(register__n1112) );
  BUFx6f_ASAP7_75t_R register___U626 ( .A(register__n6268), .Y(register__n12442) );
  BUFx4f_ASAP7_75t_R register___U627 ( .A(register__net148251), .Y(register__net64444) );
  INVx1_ASAP7_75t_R register___U628 ( .A(register__n12603), .Y(register__n93) );
  INVx2_ASAP7_75t_R register___U629 ( .A(register__n11905), .Y(register__n1524) );
  INVx4_ASAP7_75t_R register___U630 ( .A(register__n4270), .Y(register__n1549) );
  BUFx4f_ASAP7_75t_R register___U631 ( .A(register__n4270), .Y(register__n11910) );
  INVxp67_ASAP7_75t_R register___U632 ( .A(register__n4270), .Y(register__n1547) );
  BUFx4f_ASAP7_75t_R register___U633 ( .A(register__n4270), .Y(register__n1550) );
  INVx1_ASAP7_75t_R register___U634 ( .A(register__n1549), .Y(register__n734) );
  NAND2xp67_ASAP7_75t_R register___U635 ( .A(register__net64976), .B(register__n204), .Y(register__n432) );
  BUFx10_ASAP7_75t_R register___U636 ( .A(register__n11910), .Y(register__n11909) );
  INVx2_ASAP7_75t_R register___U637 ( .A(register__n1550), .Y(register__n113) );
  INVx3_ASAP7_75t_R register___U638 ( .A(register__n1962), .Y(register__n1960) );
  INVx2_ASAP7_75t_R register___U639 ( .A(register__n1517), .Y(register__n107) );
  INVx2_ASAP7_75t_R register___U640 ( .A(register__n734), .Y(register__n7088) );
  INVx1_ASAP7_75t_R register___U641 ( .A(register__n1959), .Y(register__n1535) );
  BUFx3_ASAP7_75t_R register___U642 ( .A(register__net148251), .Y(register__net144716) );
  BUFx2_ASAP7_75t_R register___U643 ( .A(register__net147584), .Y(register__net148251) );
  CKINVDCx11_ASAP7_75t_R register___U644 ( .A(register__n12066), .Y(register__n1374) );
  INVx3_ASAP7_75t_R register___U645 ( .A(register__n8561), .Y(register__n12064) );
  BUFx6f_ASAP7_75t_R register___U646 ( .A(register__n82), .Y(register__n3746) );
  BUFx12f_ASAP7_75t_R register___U647 ( .A(register__n81), .Y(register__n1992) );
  BUFx12f_ASAP7_75t_R register___U648 ( .A(register__n81), .Y(register__n3076) );
  BUFx16f_ASAP7_75t_R register___U649 ( .A(register__n3076), .Y(register__n2800) );
  CKINVDCx9p33_ASAP7_75t_R register___U650 ( .A(register__n82), .Y(register__n665) );
  CKINVDCx9p33_ASAP7_75t_R register___U651 ( .A(register__n82), .Y(register__n1069) );
  INVx4_ASAP7_75t_R register___U652 ( .A(register__n2800), .Y(register__n1946) );
  INVx2_ASAP7_75t_R register___U653 ( .A(register__n1992), .Y(register__n2801) );
  INVx4_ASAP7_75t_R register___U654 ( .A(register__n1992), .Y(register__n2799) );
  AND2x6_ASAP7_75t_R register___U655 ( .A(register__n11131), .B(register__n312), .Y(register__C6422_net59548) );
  BUFx12f_ASAP7_75t_R register___U656 ( .A(register__net130666), .Y(register__C6422_net69762) );
  BUFx4f_ASAP7_75t_R register___U657 ( .A(register__net130666), .Y(register__net109844) );
  AND2x6_ASAP7_75t_R register___U658 ( .A(register__n11135), .B(register__n312), .Y(register__C6422_net59540) );
  CKINVDCx6p67_ASAP7_75t_R register___U659 ( .A(register__net144425), .Y(register__net62678) );
  INVx6_ASAP7_75t_R register___U660 ( .A(register__net62678), .Y(register__net100799) );
  BUFx3_ASAP7_75t_R register___U661 ( .A(register__net62716), .Y(register__net141449) );
  AND2x6_ASAP7_75t_R register___U662 ( .A(register__n11141), .B(register__n312), .Y(register__C6422_net60408) );
  AND2x4_ASAP7_75t_R register___U663 ( .A(register__n12488), .B(register__n593), .Y(register__n7684) );
  AND3x4_ASAP7_75t_R register___U664 ( .A(register__n1128), .B(register__n5734), .C(register__n707), .Y(register__n12490) );
  BUFx6f_ASAP7_75t_R register___U665 ( .A(register__n3298), .Y(register__n11785) );
  BUFx5_ASAP7_75t_R register___U666 ( .A(register__n3298), .Y(register__n2829) );
  NAND2x1_ASAP7_75t_R register___U667 ( .A(register__n1963), .B(register__n12484), .Y(register__n94) );
  INVx2_ASAP7_75t_R register___U668 ( .A(register__n1563), .Y(register__n1567) );
  INVx1_ASAP7_75t_R register___U669 ( .A(register__n1563), .Y(register__n1568) );
  INVx1_ASAP7_75t_R register___U670 ( .A(register__n1563), .Y(register__n1565) );
  INVx1_ASAP7_75t_R register___U671 ( .A(register__n1563), .Y(register__n1566) );
  INVx2_ASAP7_75t_R register___U672 ( .A(register__n1563), .Y(register__n1569) );
  INVx2_ASAP7_75t_R register___U673 ( .A(register__n94), .Y(register__n1194) );
  INVx1_ASAP7_75t_R register___U674 ( .A(register__n13119), .Y(register__n95) );
  AND2x6_ASAP7_75t_R register___U675 ( .A(register__n1963), .B(register__n7684), .Y(register__n3821) );
  BUFx16f_ASAP7_75t_R register___U676 ( .A(register__n3821), .Y(register__n3336) );
  BUFx16f_ASAP7_75t_R register___U677 ( .A(register__n3821), .Y(register__n3334) );
  CKINVDCx10_ASAP7_75t_R register___U678 ( .A(register__n3335), .Y(register__n1266) );
  BUFx4f_ASAP7_75t_R register___U679 ( .A(register__n1), .Y(register__register__n11847) );
  BUFx6f_ASAP7_75t_R register___U680 ( .A(register__n12487), .Y(register__n3407) );
  INVx1_ASAP7_75t_R register___U681 ( .A(register__n12568), .Y(register__n96) );
  INVx1_ASAP7_75t_R register___U682 ( .A(register__n12569), .Y(register__n97) );
  AND2x6_ASAP7_75t_R register___U683 ( .A(register__n10518), .B(register__n12484), .Y(register__n4851) );
  XNOR2x2_ASAP7_75t_R register___U684 ( .A(register__n2277), .B(register__n1128), .Y(register__n12505) );
  AND3x2_ASAP7_75t_R register___U685 ( .A(register__n5301), .B(register__n707), .C(register__n12488), .Y(register__n796) );
  OR3x2_ASAP7_75t_R register___U686 ( .A(WB_rd[0]), .B(WB_rd[2]), .C(
        WB_rd[1]), .Y(register__n12491) );
  INVx1_ASAP7_75t_R register___U687 ( .A(register__n600), .Y(register__n98) );
  INVx2_ASAP7_75t_R register___U688 ( .A(register__n3706), .Y(register__n600) );
  AND3x2_ASAP7_75t_R register___U689 ( .A(register__n5301), .B(register__n12489), .C(WB_rd[0]), .Y(
        n12487) );
  INVx2_ASAP7_75t_R register___U690 ( .A(register__n7327), .Y(register__n1306) );
  INVx4_ASAP7_75t_R register___U691 ( .A(register__n7327), .Y(register__n598) );
  CKINVDCx6p67_ASAP7_75t_R register___U692 ( .A(WB_rd[2]), .Y(register__n707) );
  AND3x4_ASAP7_75t_R register___U693 ( .A(register__n5049), .B(register__n12502), .C(register__n666), .Y(register__n12503) );
  NAND3x2_ASAP7_75t_R register___U694 ( .A(WB_rd[1]), .B(register__n707), .C(register__n12488), .Y(
        n1503) );
  INVx6_ASAP7_75t_R register___U695 ( .A(register__n5173), .Y(register__n1120) );
  NOR2x1p5_ASAP7_75t_R register___U696 ( .A(register__n1036), .B(register__n11727), .Y(register__n1074) );
  INVx4_ASAP7_75t_R register___U697 ( .A(register__n5548), .Y(register__n1792) );
  AND2x6_ASAP7_75t_R register___U698 ( .A(register__n385), .B(register__n12490), .Y(register__n5548) );
  INVx3_ASAP7_75t_R register___U699 ( .A(register__n12336), .Y(register__n12322) );
  INVx4_ASAP7_75t_R register___U700 ( .A(register__n5351), .Y(register__n12336) );
  INVx3_ASAP7_75t_R register___U701 ( .A(register__net62684), .Y(register__net62660) );
  BUFx12f_ASAP7_75t_R register___U702 ( .A(register__net62718), .Y(register__net62684) );
  AND2x6_ASAP7_75t_R register___U703 ( .A(register__n6467), .B(register__n12503), .Y(register__n12504) );
  INVx1_ASAP7_75t_R register___U704 ( .A(register__n5550), .Y(register__n1740) );
  INVx1_ASAP7_75t_R register___U705 ( .A(register__n5878), .Y(register__n1427) );
  INVx1_ASAP7_75t_R register___U706 ( .A(register__n5650), .Y(register__n1393) );
  INVx1_ASAP7_75t_R register___U707 ( .A(register__n5208), .Y(register__n1264) );
  INVx3_ASAP7_75t_R register___U708 ( .A(register__n5185), .Y(register__n99) );
  BUFx8_ASAP7_75t_R register___U709 ( .A(register__n1746), .Y(register__n100) );
  BUFx8_ASAP7_75t_R register___U710 ( .A(register__n1747), .Y(register__n101) );
  INVx3_ASAP7_75t_R register___U711 ( .A(register__n2115), .Y(register__n2116) );
  BUFx10_ASAP7_75t_R register___U712 ( .A(register__n12493), .Y(register__n1138) );
  CKINVDCx10_ASAP7_75t_R register___U713 ( .A(register__n1138), .Y(register__n103) );
  INVx1_ASAP7_75t_R register___U714 ( .A(register__n1413), .Y(register__n1333) );
  INVx3_ASAP7_75t_R register___U715 ( .A(register__n5548), .Y(register__n1794) );
  INVx4_ASAP7_75t_R register___U716 ( .A(register__n5548), .Y(register__n11815) );
  INVx3_ASAP7_75t_R register___U717 ( .A(register__n5548), .Y(register__n1643) );
  INVx3_ASAP7_75t_R register___U718 ( .A(register__n1625), .Y(register__n104) );
  INVx5_ASAP7_75t_R register___U719 ( .A(register__n11814), .Y(register__n1625) );
  HB1xp67_ASAP7_75t_R register___U720 ( .A(register__n2119), .Y(register__n105) );
  HB1xp67_ASAP7_75t_R register___U721 ( .A(register__n2119), .Y(register__n106) );
  BUFx10_ASAP7_75t_R register___U722 ( .A(register__n3376), .Y(register__n108) );
  BUFx2_ASAP7_75t_R register___U723 ( .A(register__n12184), .Y(register__n3376) );
  BUFx16f_ASAP7_75t_R register___U724 ( .A(register__n3021), .Y(register__n1583) );
  CKINVDCx20_ASAP7_75t_R register___U725 ( .A(register__n1583), .Y(register__n109) );
  INVx5_ASAP7_75t_R register___U726 ( .A(register__n1664), .Y(register__n114) );
  INVx2_ASAP7_75t_R register___U727 ( .A(register__net146710), .Y(register__n1664) );
  INVx5_ASAP7_75t_R register___U728 ( .A(register__n1624), .Y(register__n115) );
  INVx2_ASAP7_75t_R register___U729 ( .A(register__n11893), .Y(register__n1624) );
  CKINVDCx5p33_ASAP7_75t_R register___U730 ( .A(register__n1654), .Y(register__n116) );
  BUFx4_ASAP7_75t_R register___U731 ( .A(register__n94), .Y(register__n118) );
  BUFx2_ASAP7_75t_R register___U732 ( .A(register__net94610), .Y(register__net113148) );
  BUFx4_ASAP7_75t_R register___U733 ( .A(register__n1547), .Y(register__n119) );
  BUFx12_ASAP7_75t_R register___U734 ( .A(register__n1567), .Y(register__n120) );
  BUFx3_ASAP7_75t_R register___U735 ( .A(register__n7996), .Y(register__n441) );
  INVx1_ASAP7_75t_R register___U736 ( .A(register__net109611), .Y(register__n1986) );
  NAND2xp5_ASAP7_75t_R register___U737 ( .A(register__net123879), .B(register__net89421), .Y(register__n2678) );
  OAI22xp33_ASAP7_75t_R register___U738 ( .A1(register__register__n12148), .A2(register__n1549), .B1(register__n9752), .B2(register__n1532), 
        .Y(register__n121) );
  BUFx6f_ASAP7_75t_R register___U739 ( .A(register__n3604), .Y(register__n3514) );
  HB1xp67_ASAP7_75t_R register___U740 ( .A(register__n13079), .Y(register__n4891) );
  NOR2xp67_ASAP7_75t_R register___U741 ( .A(register__n2278), .B(register__n2279), .Y(register__n122) );
  NOR3xp33_ASAP7_75t_R register___U742 ( .A(register__n123), .B(register__n11322), .C(register__n2280), .Y(register__n6161) );
  INVxp67_ASAP7_75t_R register___U743 ( .A(register__n122), .Y(register__n123) );
  INVx1_ASAP7_75t_R register___U744 ( .A(register__n11321), .Y(register__n2279) );
  INVx1_ASAP7_75t_R register___U745 ( .A(register__n11320), .Y(register__n2278) );
  NOR2x1_ASAP7_75t_R register___U746 ( .A(register__n1278), .B(register__n1304), .Y(register__n7614) );
  CKINVDCx6p67_ASAP7_75t_R register___U747 ( .A(register__n514), .Y(register__n515) );
  INVx5_ASAP7_75t_R register___U748 ( .A(register__net94400), .Y(register__n514) );
  HB1xp67_ASAP7_75t_R register___U749 ( .A(register__n11388), .Y(register__n5818) );
  HB1xp67_ASAP7_75t_R register___U750 ( .A(register__n11323), .Y(register__n5327) );
  INVx1_ASAP7_75t_R register___U751 ( .A(register__n5298), .Y(register__n124) );
  AO22x1_ASAP7_75t_R register___U752 ( .A1(register__net90665), .A2(register__net91683), .B1(register__net89617), .B2(
        n1352), .Y(register__n10724) );
  AO22x1_ASAP7_75t_R register___U753 ( .A1(register__n9409), .A2(register__net91683), .B1(register__net96692), .B2(
        n9423), .Y(register__n10830) );
  AO22x1_ASAP7_75t_R register___U754 ( .A1(register__n1249), .A2(register__n4579), .B1(register__n125), .B2(register__n1120), .Y(
        n383) );
  CKINVDCx20_ASAP7_75t_R register___U755 ( .A(register__n9867), .Y(register__n125) );
  INVxp67_ASAP7_75t_R register___U756 ( .A(register__n1249), .Y(register__n12398) );
  INVx1_ASAP7_75t_R register___U757 ( .A(register__n10998), .Y(register__n126) );
  HB1xp67_ASAP7_75t_R register___U758 ( .A(register__n12484), .Y(register__n3940) );
  OR2x2_ASAP7_75t_R register___U759 ( .A(register__n1036), .B(register__n7697), .Y(register__n127) );
  BUFx6f_ASAP7_75t_R register___U760 ( .A(register__n268), .Y(register__n128) );
  OR2x2_ASAP7_75t_R register___U761 ( .A(register__n653), .B(register__n7697), .Y(register__n129) );
  BUFx6f_ASAP7_75t_R register___U762 ( .A(register__n12497), .Y(register__n3298) );
  INVxp67_ASAP7_75t_R register___U763 ( .A(register__n12497), .Y(register__n1576) );
  OAI22xp5_ASAP7_75t_R register___U764 ( .A1(register__n1949), .A2(register__n3721), .B1(register__n6059), .B2(register__n1687), 
        .Y(read_reg_data_2[28]) );
  HB1xp67_ASAP7_75t_R register___U765 ( .A(register__n3294), .Y(register__n3293) );
  INVx1_ASAP7_75t_R register___U766 ( .A(register__register__n13089), .Y(register__n130) );
  OAI22xp33_ASAP7_75t_R register___U767 ( .A1(register__n12148), .A2(register__n3991), .B1(register__n6096), .B2(register__n4843), 
        .Y(register__n131) );
  INVx4_ASAP7_75t_R register___U768 ( .A(register__net62684), .Y(register__net119634) );
  INVx5_ASAP7_75t_R register___U769 ( .A(register__net119634), .Y(register__net125327) );
  BUFx3_ASAP7_75t_R register___U770 ( .A(register__n883), .Y(register__net125426) );
  INVx2_ASAP7_75t_R register___U771 ( .A(register__n3205), .Y(register__n7908) );
  OAI22xp33_ASAP7_75t_R register___U772 ( .A1(register__net66310), .A2(register__n9176), .B1(register__n12206), .B2(
        n1687), .Y(read_reg_data_2[16]) );
  INVxp67_ASAP7_75t_R register___U773 ( .A(register__n7697), .Y(register__n772) );
  OR2x2_ASAP7_75t_R register___U774 ( .A(register__n1335), .B(register__n7697), .Y(register__n275) );
  BUFx4f_ASAP7_75t_R register___U775 ( .A(register__n12109), .Y(register__n4004) );
  BUFx6f_ASAP7_75t_R register___U776 ( .A(register__n12109), .Y(register__n5034) );
  INVx3_ASAP7_75t_R register___U777 ( .A(write_data[9]), .Y(register__n12109) );
  AO22x1_ASAP7_75t_R register___U778 ( .A1(register__net62682), .A2(register__n4851), .B1(register__n133), .B2(register__n809), 
        .Y(register__n132) );
  CKINVDCx20_ASAP7_75t_R register___U779 ( .A(register__n10417), .Y(register__n133) );
  INVx1_ASAP7_75t_R register___U780 ( .A(register__n4851), .Y(register__n701) );
  HB1xp67_ASAP7_75t_R register___U781 ( .A(register__n9065), .Y(register__n6044) );
  BUFx6f_ASAP7_75t_R register___U782 ( .A(register__n5524), .Y(register__n11831) );
  INVxp67_ASAP7_75t_R register___U783 ( .A(register__n11143), .Y(register__n572) );
  HB1xp67_ASAP7_75t_R register___U784 ( .A(register__n11186), .Y(register__n4735) );
  AO22x1_ASAP7_75t_R register___U785 ( .A1(register__net90253), .A2(register__C6423_net61318), .B1(register__net100896), 
        .B2(register__n1449), .Y(register__n11608) );
  AO22x1_ASAP7_75t_R register___U786 ( .A1(register__n9256), .A2(register__C6423_net61318), .B1(register__n10028), .B2(
        n1449), .Y(register__n11209) );
  BUFx10_ASAP7_75t_R register___U787 ( .A(register__net146267), .Y(register__net64456) );
  OAI22xp33_ASAP7_75t_R register___U788 ( .A1(register__n12148), .A2(register__n951), .B1(register__n958), .B2(register__n9744), 
        .Y(register__n134) );
  INVx1_ASAP7_75t_R register___U789 ( .A(register__n12801), .Y(register__n135) );
  BUFx2_ASAP7_75t_R register___U790 ( .A(register__n12250), .Y(register__n4290) );
  INVx2_ASAP7_75t_R register___U791 ( .A(write_data[7]), .Y(register__net144804) );
  AND2x6_ASAP7_75t_R register___U792 ( .A(register__n312), .B(register__n612), .Y(register__n1771) );
  NOR2xp33_ASAP7_75t_R register___U793 ( .A(register__n1803), .B(register__n1802), .Y(register__n136) );
  NOR2xp33_ASAP7_75t_R register___U794 ( .A(register__n1801), .B(register__n137), .Y(register__n5318) );
  INVxp33_ASAP7_75t_R register___U795 ( .A(register__n136), .Y(register__n137) );
  NOR2xp33_ASAP7_75t_R register___U796 ( .A(register__n1987), .B(register__n10958), .Y(register__n1801) );
  NOR2xp33_ASAP7_75t_R register___U797 ( .A(register__n1995), .B(register__n10959), .Y(register__n1802) );
  NOR2xp33_ASAP7_75t_R register___U798 ( .A(register__n1800), .B(register__n10960), .Y(register__n1803) );
  INVx1_ASAP7_75t_R register___U799 ( .A(register__n1833), .Y(register__n1834) );
  INVx1_ASAP7_75t_R register___U800 ( .A(register__n13320), .Y(register__n138) );
  NOR2xp33_ASAP7_75t_R register___U801 ( .A(register__n420), .B(register__n8836), .Y(register__n797) );
  CKINVDCx10_ASAP7_75t_R register___U802 ( .A(register__n11998), .Y(register__n6405) );
  HB1xp67_ASAP7_75t_R register___U803 ( .A(register__n12885), .Y(register__n4057) );
  INVx1_ASAP7_75t_R register___U804 ( .A(register__n127), .Y(register__n284) );
  BUFx4f_ASAP7_75t_R register___U805 ( .A(register__net122862), .Y(register__C6423_net68766) );
  HB1xp67_ASAP7_75t_R register___U806 ( .A(register__n3163), .Y(register__n3162) );
  INVx2_ASAP7_75t_R register___U807 ( .A(register__n1958), .Y(register__n1959) );
  INVxp67_ASAP7_75t_R register___U808 ( .A(register__n11356), .Y(register__n5744) );
  HB1xp67_ASAP7_75t_R register___U809 ( .A(register__net94400), .Y(register__n235) );
  HB1xp67_ASAP7_75t_R register___U810 ( .A(register__n6270), .Y(register__n6758) );
  INVx1_ASAP7_75t_R register___U811 ( .A(register__n13142), .Y(register__n140) );
  INVxp33_ASAP7_75t_R register___U812 ( .A(register__net150703), .Y(register__n157) );
  INVx3_ASAP7_75t_R register___U813 ( .A(register__n277), .Y(register__n1999) );
  BUFx4f_ASAP7_75t_R register___U814 ( .A(register__n277), .Y(register__net104679) );
  BUFx2_ASAP7_75t_R register___U815 ( .A(register__n2894), .Y(register__n2893) );
  BUFx3_ASAP7_75t_R register___U816 ( .A(register__n5227), .Y(register__n5226) );
  BUFx2_ASAP7_75t_R register___U817 ( .A(register__n5227), .Y(register__n3842) );
  INVx2_ASAP7_75t_R register___U818 ( .A(register__n3348), .Y(register__n245) );
  NAND2xp67_ASAP7_75t_R register___U819 ( .A(register__n3348), .B(register__n3344), .Y(register__n1154) );
  BUFx4f_ASAP7_75t_R register___U820 ( .A(write_data[20]), .Y(register__n5351) );
  INVx6_ASAP7_75t_R register___U821 ( .A(register__n5497), .Y(register__n12315) );
  BUFx12f_ASAP7_75t_R register___U822 ( .A(register__n3572), .Y(register__n3258) );
  BUFx5_ASAP7_75t_R register___U823 ( .A(register__C6423_net61343), .Y(register__net122249) );
  NOR2xp67_ASAP7_75t_R register___U824 ( .A(register__n10817), .B(register__n142), .Y(register__n1744) );
  NAND2xp67_ASAP7_75t_R register___U825 ( .A(register__n2788), .B(register__n1745), .Y(register__n142) );
  BUFx2_ASAP7_75t_R register___U826 ( .A(register__n1161), .Y(register__n5343) );
  BUFx2_ASAP7_75t_R register___U827 ( .A(register__n1161), .Y(register__n3651) );
  BUFx2_ASAP7_75t_R register___U828 ( .A(register__n1161), .Y(register__n3680) );
  BUFx3_ASAP7_75t_R register___U829 ( .A(register__n1161), .Y(register__n5341) );
  INVx5_ASAP7_75t_R register___U830 ( .A(register__n3336), .Y(register__n1755) );
  BUFx2_ASAP7_75t_R register___U831 ( .A(register__n732), .Y(register__n12248) );
  BUFx5_ASAP7_75t_R register___U832 ( .A(register__n3571), .Y(register__n3474) );
  INVx1_ASAP7_75t_R register___U833 ( .A(register__n12963), .Y(register__n143) );
  INVx3_ASAP7_75t_R register___U834 ( .A(write_data[16]), .Y(register__n12224) );
  OAI22xp33_ASAP7_75t_R register___U835 ( .A1(register__n12456), .A2(register__n1092), .B1(register__n9756), .B2(register__n5530), 
        .Y(register__n144) );
  INVxp33_ASAP7_75t_R register___U836 ( .A(register__n11943), .Y(register__n145) );
  BUFx3_ASAP7_75t_R register___U837 ( .A(register__n11948), .Y(register__n4377) );
  BUFx2_ASAP7_75t_R register___U838 ( .A(register__n11941), .Y(register__n11943) );
  INVx2_ASAP7_75t_R register___U839 ( .A(register__C6423_net61355), .Y(register__net150876) );
  NOR2xp33_ASAP7_75t_R register___U840 ( .A(register__net62664), .B(register__n1974), .Y(register__n146) );
  NOR2xp33_ASAP7_75t_R register___U841 ( .A(register__n10467), .B(register__n2843), .Y(register__n147) );
  NOR2xp33_ASAP7_75t_R register___U842 ( .A(register__n146), .B(register__n147), .Y(register__n12888) );
  INVxp67_ASAP7_75t_R register___U843 ( .A(register__n12888), .Y(register__n148) );
  INVxp67_ASAP7_75t_R register___U844 ( .A(register__n11143), .Y(register__n565) );
  INVx1_ASAP7_75t_R register___U845 ( .A(register__n7697), .Y(register__n8337) );
  NOR2xp33_ASAP7_75t_R register___U846 ( .A(register__n2003), .B(register__n2611), .Y(register__n2612) );
  INVxp33_ASAP7_75t_R register___U847 ( .A(register__n2003), .Y(register__net150894) );
  INVx1_ASAP7_75t_R register___U848 ( .A(register__n1998), .Y(register__n2003) );
  HB1xp67_ASAP7_75t_R register___U849 ( .A(register__n12829), .Y(register__n3766) );
  CKINVDCx10_ASAP7_75t_R register___U850 ( .A(register__n4199), .Y(register__n11998) );
  INVx2_ASAP7_75t_R register___U851 ( .A(rs2[3]), .Y(register__n1432) );
  AND2x2_ASAP7_75t_R register___U852 ( .A(register__n5441), .B(register__n2744), .Y(register__n149) );
  AND2x2_ASAP7_75t_R register___U853 ( .A(register__n5441), .B(register__n2744), .Y(register__n740) );
  BUFx2_ASAP7_75t_R register___U854 ( .A(register__n5443), .Y(register__n3364) );
  BUFx3_ASAP7_75t_R register___U855 ( .A(register__n12224), .Y(register__n5443) );
  NOR2x1_ASAP7_75t_R register___U856 ( .A(register__n2780), .B(register__n2781), .Y(register__n12739) );
  INVx1_ASAP7_75t_R register___U857 ( .A(register__n12739), .Y(register__n2249) );
  AND2x6_ASAP7_75t_R register___U858 ( .A(register__n1107), .B(register__n11728), .Y(register__net110414) );
  INVx1_ASAP7_75t_R register___U859 ( .A(n9), .Y(register__n12250) );
  NAND2xp33_ASAP7_75t_R register___U860 ( .A(register__n6966), .B(register__net122579), .Y(register__n150) );
  NAND2xp33_ASAP7_75t_R register___U861 ( .A(register__n10289), .B(register__n1998), .Y(register__n151) );
  NAND2xp33_ASAP7_75t_R register___U862 ( .A(register__n150), .B(register__n151), .Y(register__n11635) );
  HB1xp67_ASAP7_75t_R register___U863 ( .A(register__n9311), .Y(register__n6966) );
  BUFx6f_ASAP7_75t_R register___U864 ( .A(register__n9099), .Y(register__n10289) );
  INVx1_ASAP7_75t_R register___U865 ( .A(register__n11360), .Y(register__n152) );
  NAND2x1p5_ASAP7_75t_R register___U866 ( .A(rs2[4]), .B(register__n1432), .Y(register__n653) );
  AND2x6_ASAP7_75t_R register___U867 ( .A(register__n1953), .B(register__n11719), .Y(register__net125170) );
  NOR3xp33_ASAP7_75t_R register___U868 ( .A(register__n30), .B(register__n2357), .C(register__n2368), .Y(register__n2319) );
  NOR2xp33_ASAP7_75t_R register___U869 ( .A(register__net126596), .B(register__n2329), .Y(register__n2330) );
  BUFx2_ASAP7_75t_R register___U870 ( .A(register__n4121), .Y(register__n4120) );
  NOR2xp67_ASAP7_75t_R register___U871 ( .A(register__net150876), .B(register__n2434), .Y(register__n2435) );
  INVxp33_ASAP7_75t_R register___U872 ( .A(register__net150876), .Y(register__net150888) );
  INVxp67_ASAP7_75t_R register___U873 ( .A(register__n1432), .Y(register__n821) );
  BUFx2_ASAP7_75t_R register___U874 ( .A(register__n821), .Y(register__n1011) );
  INVx1_ASAP7_75t_R register___U875 ( .A(register__n1687), .Y(register__n1553) );
  BUFx16f_ASAP7_75t_R register___U876 ( .A(register__net61445), .Y(register__n1687) );
  AND2x6_ASAP7_75t_R register___U877 ( .A(register__n1552), .B(register__n1553), .Y(register__n1251) );
  BUFx6f_ASAP7_75t_R register___U878 ( .A(register__net64444), .Y(register__net146408) );
  HB1xp67_ASAP7_75t_R register___U879 ( .A(register__n10810), .Y(register__n4166) );
  INVxp67_ASAP7_75t_R register___U880 ( .A(register__n11635), .Y(register__n6425) );
  OR2x2_ASAP7_75t_R register___U881 ( .A(register__n653), .B(register__n7697), .Y(register__n153) );
  OR2x2_ASAP7_75t_R register___U882 ( .A(register__n653), .B(register__n7697), .Y(register__n762) );
  AOI222xp33_ASAP7_75t_R register___U883 ( .A1(register__net109611), .A2(register__n10347), .B1(register__n1993), .B2(
        n9439), .C1(register__n831), .C2(register__n7127), .Y(register__n11323) );
  INVx5_ASAP7_75t_R register___U884 ( .A(register__n1800), .Y(register__n831) );
  INVx2_ASAP7_75t_R register___U885 ( .A(register__n10665), .Y(register__n9156) );
  BUFx4_ASAP7_75t_R register___U886 ( .A(register__n7128), .Y(register__n7127) );
  INVxp67_ASAP7_75t_R register___U887 ( .A(register__n507), .Y(register__n155) );
  INVxp33_ASAP7_75t_R register___U888 ( .A(register__n37), .Y(register__net150703) );
  AND2x4_ASAP7_75t_R register___U889 ( .A(register__n12490), .B(register__n1985), .Y(register__n7050) );
  BUFx4f_ASAP7_75t_R register___U890 ( .A(register__n6268), .Y(register__n12449) );
  INVx2_ASAP7_75t_R register___U891 ( .A(register__n5286), .Y(register__n7638) );
  BUFx6f_ASAP7_75t_R register___U892 ( .A(register__net116957), .Y(register__net66302) );
  HB1xp67_ASAP7_75t_R register___U893 ( .A(Reg_data[349]), .Y(register__net94810) );
  INVx1_ASAP7_75t_R register___U894 ( .A(register__n11081), .Y(register__n8295) );
  HB1xp67_ASAP7_75t_R register___U895 ( .A(register__n11948), .Y(register__n4816) );
  BUFx12f_ASAP7_75t_R register___U896 ( .A(register__n3538), .Y(register__n3536) );
  BUFx4f_ASAP7_75t_R register___U897 ( .A(register__n3842), .Y(register__n5224) );
  BUFx6f_ASAP7_75t_R register___U898 ( .A(register__n12495), .Y(register__n385) );
  INVx2_ASAP7_75t_R register___U899 ( .A(register__n1981), .Y(register__n1958) );
  INVx1_ASAP7_75t_R register___U900 ( .A(register__C6423_net60460), .Y(register__n712) );
  NOR2x1_ASAP7_75t_R register___U901 ( .A(register__n5441), .B(register__n1133), .Y(register__n883) );
  INVx1_ASAP7_75t_R register___U902 ( .A(register__n1345), .Y(register__n1353) );
  BUFx3_ASAP7_75t_R register___U903 ( .A(register__n11141), .Y(register__n655) );
  HB1xp67_ASAP7_75t_R register___U904 ( .A(register__n12534), .Y(register__n4217) );
  INVx2_ASAP7_75t_R register___U905 ( .A(register__n2015), .Y(register__n1113) );
  INVx2_ASAP7_75t_R register___U906 ( .A(register__n2015), .Y(register__net149934) );
  INVx2_ASAP7_75t_R register___U907 ( .A(register__n2015), .Y(register__net149937) );
  INVx1_ASAP7_75t_R register___U908 ( .A(register__n2015), .Y(register__n1114) );
  INVxp67_ASAP7_75t_R register___U909 ( .A(register__n5128), .Y(register__n8305) );
  CKINVDCx5p33_ASAP7_75t_R register___U910 ( .A(register__n488), .Y(register__C6423_net61335) );
  BUFx3_ASAP7_75t_R register___U911 ( .A(register__n5514), .Y(register__n4282) );
  HB1xp67_ASAP7_75t_R register___U912 ( .A(register__n3948), .Y(register__n5514) );
  INVx3_ASAP7_75t_R register___U913 ( .A(register__n3948), .Y(register__n12254) );
  BUFx2_ASAP7_75t_R register___U914 ( .A(register__n12277), .Y(register__n3948) );
  INVx1_ASAP7_75t_R register___U915 ( .A(register__n13340), .Y(register__n160) );
  HB1xp67_ASAP7_75t_R register___U916 ( .A(register__n5600), .Y(register__n5599) );
  HB1xp67_ASAP7_75t_R register___U917 ( .A(register__n5784), .Y(register__n5783) );
  INVxp67_ASAP7_75t_R register___U918 ( .A(register__n7354), .Y(register__n8597) );
  HB1xp67_ASAP7_75t_R register___U919 ( .A(register__n7355), .Y(register__n7354) );
  OAI22xp33_ASAP7_75t_R register___U920 ( .A1(register__n12433), .A2(register__n4267), .B1(register__n9897), .B2(register__n4841), 
        .Y(register__n161) );
  NOR2xp67_ASAP7_75t_R register___U921 ( .A(register__n11221), .B(register__n279), .Y(register__n278) );
  INVx1_ASAP7_75t_R register___U922 ( .A(register__n262), .Y(register__n263) );
  CKINVDCx12_ASAP7_75t_R register___U923 ( .A(register__n1771), .Y(register__n1558) );
  HB1xp67_ASAP7_75t_R register___U924 ( .A(register__net122862), .Y(register__n162) );
  BUFx2_ASAP7_75t_R register___U925 ( .A(register__net125804), .Y(register__C6423_net68764) );
  BUFx6f_ASAP7_75t_R register___U926 ( .A(register__C6423_net68766), .Y(register__net125803) );
  BUFx2_ASAP7_75t_R register___U927 ( .A(register__net139882), .Y(register__net139058) );
  INVx1_ASAP7_75t_R register___U928 ( .A(register__C6422_net60443), .Y(register__n367) );
  NOR2xp67_ASAP7_75t_R register___U929 ( .A(register__net64350), .B(register__n399), .Y(register__n615) );
  NOR2xp67_ASAP7_75t_R register___U930 ( .A(register__n615), .B(register__n616), .Y(register__n13300) );
  BUFx3_ASAP7_75t_R register___U931 ( .A(register__net64398), .Y(register__net147144) );
  INVx1_ASAP7_75t_R register___U932 ( .A(register__n12968), .Y(register__n163) );
  BUFx6f_ASAP7_75t_R register___U933 ( .A(register__n3915), .Y(register__n12301) );
  INVx1_ASAP7_75t_R register___U934 ( .A(register__n12563), .Y(register__n164) );
  INVx1_ASAP7_75t_R register___U935 ( .A(register__n12218), .Y(register__n12202) );
  INVx4_ASAP7_75t_R register___U936 ( .A(register__n3729), .Y(register__n12432) );
  INVx2_ASAP7_75t_R register___U937 ( .A(register__n2167), .Y(register__n10518) );
  INVxp67_ASAP7_75t_R register___U938 ( .A(register__n3026), .Y(register__n4486) );
  NAND2xp67_ASAP7_75t_R register___U939 ( .A(register__n518), .B(register__n2412), .Y(read_reg_data_2[25]) );
  AO22x1_ASAP7_75t_R register___U940 ( .A1(register__n9648), .A2(register__n3), .B1(register__n9975), .B2(register__n233), .Y(
        n10677) );
  OAI22xp33_ASAP7_75t_R register___U941 ( .A1(register__n12376), .A2(register__n698), .B1(register__n9487), .B2(register__n688), 
        .Y(register__n165) );
  INVx3_ASAP7_75t_R register___U942 ( .A(register__C6423_net60462), .Y(register__n353) );
  INVx1_ASAP7_75t_R register___U943 ( .A(register__n13209), .Y(register__n166) );
  INVx2_ASAP7_75t_R register___U944 ( .A(register__n11945), .Y(register__n11933) );
  BUFx2_ASAP7_75t_R register___U945 ( .A(register__n5443), .Y(register__n12217) );
  BUFx4f_ASAP7_75t_R register___U946 ( .A(register__n5443), .Y(register__n3320) );
  INVxp67_ASAP7_75t_R register___U947 ( .A(register__n4218), .Y(register__n6445) );
  OAI22xp33_ASAP7_75t_R register___U948 ( .A1(register__n145), .A2(register__n3719), .B1(register__n10363), .B2(register__n1164), 
        .Y(register__n167) );
  BUFx4f_ASAP7_75t_R register___U949 ( .A(register__n3602), .Y(register__n3915) );
  BUFx6f_ASAP7_75t_R register___U950 ( .A(register__n3602), .Y(register__n12308) );
  INVx2_ASAP7_75t_R register___U951 ( .A(register__n4015), .Y(register__n6406) );
  BUFx6f_ASAP7_75t_R register___U952 ( .A(register__n3538), .Y(register__n3537) );
  HB1xp67_ASAP7_75t_R register___U953 ( .A(register__n1226), .Y(register__n168) );
  INVxp33_ASAP7_75t_R register___U954 ( .A(register__n1226), .Y(register__n169) );
  HB1xp67_ASAP7_75t_R register___U955 ( .A(register__n1226), .Y(register__net134749) );
  OAI22xp33_ASAP7_75t_R register___U956 ( .A1(register__n12433), .A2(register__n114), .B1(register__n10419), .B2(register__n1664), 
        .Y(register__n170) );
  BUFx6f_ASAP7_75t_R register___U957 ( .A(register__n4816), .Y(register__n11945) );
  AND3x1_ASAP7_75t_R register___U958 ( .A(register__n172), .B(register__n5138), .C(register__n10759), .Y(register__n171) );
  OA222x2_ASAP7_75t_R register___U959 ( .A1(register__n2002), .A2(register__n6220), .B1(register__n1997), .B2(register__n9158), 
        .C1(register__C6422_net69812), .C2(register__n7089), .Y(register__n172) );
  INVx6_ASAP7_75t_R register___U960 ( .A(register__n4000), .Y(register__n12461) );
  INVxp33_ASAP7_75t_R register___U961 ( .A(register__n6465), .Y(register__n1529) );
  INVx4_ASAP7_75t_R register___U962 ( .A(register__n6465), .Y(register__n11825) );
  AOI21xp5_ASAP7_75t_R register___U963 ( .A1(register__C6423_net69198), .A2(register__net90061), .B(register__n2452), 
        .Y(register__n2451) );
  NAND2xp5_ASAP7_75t_R register___U964 ( .A(register__n1744), .B(register__n2755), .Y(register__n1742) );
  AND2x2_ASAP7_75t_R register___U965 ( .A(register__n437), .B(register__n11135), .Y(register__C6422_net59544) );
  HB1xp67_ASAP7_75t_R register___U966 ( .A(Reg_data[577]), .Y(register__n6270) );
  BUFx6f_ASAP7_75t_R register___U967 ( .A(register__n3375), .Y(register__n5043) );
  OAI22xp33_ASAP7_75t_R register___U968 ( .A1(register__n12288), .A2(register__n109), .B1(register__n10112), .B2(register__n3546), 
        .Y(register__n173) );
  BUFx2_ASAP7_75t_R register___U969 ( .A(IF_ID_rs1[2]), .Y(register__n1422) );
  INVx1_ASAP7_75t_R register___U970 ( .A(register__n1111), .Y(register__n174) );
  INVxp67_ASAP7_75t_R register___U971 ( .A(register__n174), .Y(register__n175) );
  INVxp67_ASAP7_75t_R register___U972 ( .A(register__n174), .Y(register__n176) );
  INVxp67_ASAP7_75t_R register___U973 ( .A(register__n174), .Y(register__n177) );
  INVxp67_ASAP7_75t_R register___U974 ( .A(register__n174), .Y(register__n178) );
  INVxp67_ASAP7_75t_R register___U975 ( .A(register__n174), .Y(register__n179) );
  INVx1_ASAP7_75t_R register___U976 ( .A(register__n11898), .Y(register__n180) );
  INVxp67_ASAP7_75t_R register___U977 ( .A(register__n180), .Y(register__n181) );
  INVxp67_ASAP7_75t_R register___U978 ( .A(register__n180), .Y(register__n182) );
  INVxp33_ASAP7_75t_R register___U979 ( .A(register__n180), .Y(register__n183) );
  INVxp33_ASAP7_75t_R register___U980 ( .A(register__n180), .Y(register__n184) );
  INVxp33_ASAP7_75t_R register___U981 ( .A(register__n180), .Y(register__n185) );
  CKINVDCx11_ASAP7_75t_R register___U982 ( .A(register__n11896), .Y(register__n186) );
  INVx2_ASAP7_75t_R register___U983 ( .A(register__n186), .Y(register__n187) );
  INVx2_ASAP7_75t_R register___U984 ( .A(register__n186), .Y(register__n188) );
  INVx2_ASAP7_75t_R register___U985 ( .A(register__n186), .Y(register__n189) );
  INVx2_ASAP7_75t_R register___U986 ( .A(register__n186), .Y(register__n190) );
  INVx2_ASAP7_75t_R register___U987 ( .A(register__n186), .Y(register__n191) );
  INVx6_ASAP7_75t_R register___U988 ( .A(register__n3151), .Y(register__n192) );
  INVx1_ASAP7_75t_R register___U989 ( .A(register__n192), .Y(register__n193) );
  INVx1_ASAP7_75t_R register___U990 ( .A(register__n192), .Y(register__n194) );
  INVxp67_ASAP7_75t_R register___U991 ( .A(register__n192), .Y(register__n195) );
  INVx1_ASAP7_75t_R register___U992 ( .A(register__n192), .Y(register__n196) );
  INVx2_ASAP7_75t_R register___U993 ( .A(register__n192), .Y(register__n197) );
  INVxp33_ASAP7_75t_R register___U994 ( .A(register__n6302), .Y(register__n198) );
  INVxp33_ASAP7_75t_R register___U995 ( .A(register__n6302), .Y(register__n199) );
  INVxp33_ASAP7_75t_R register___U996 ( .A(register__n6302), .Y(register__n200) );
  INVxp33_ASAP7_75t_R register___U997 ( .A(register__n6302), .Y(register__n201) );
  INVxp33_ASAP7_75t_R register___U998 ( .A(register__n6302), .Y(register__n202) );
  INVxp33_ASAP7_75t_R register___U999 ( .A(register__n6302), .Y(register__n203) );
  INVxp33_ASAP7_75t_R register___U1000 ( .A(register__n198), .Y(register__n204) );
  INVxp33_ASAP7_75t_R register___U1001 ( .A(register__n198), .Y(register__n205) );
  INVxp33_ASAP7_75t_R register___U1002 ( .A(register__n198), .Y(register__n206) );
  INVxp33_ASAP7_75t_R register___U1003 ( .A(register__n199), .Y(register__n207) );
  INVxp33_ASAP7_75t_R register___U1004 ( .A(register__n199), .Y(register__n208) );
  INVxp33_ASAP7_75t_R register___U1005 ( .A(register__n199), .Y(register__n209) );
  INVxp33_ASAP7_75t_R register___U1006 ( .A(register__n200), .Y(register__n210) );
  INVxp33_ASAP7_75t_R register___U1007 ( .A(register__n200), .Y(register__n211) );
  INVxp33_ASAP7_75t_R register___U1008 ( .A(register__n200), .Y(register__n212) );
  INVxp33_ASAP7_75t_R register___U1009 ( .A(register__n201), .Y(register__n213) );
  INVxp33_ASAP7_75t_R register___U1010 ( .A(register__n201), .Y(register__n214) );
  INVxp33_ASAP7_75t_R register___U1011 ( .A(register__n201), .Y(register__n215) );
  INVxp33_ASAP7_75t_R register___U1012 ( .A(register__n202), .Y(register__n216) );
  INVxp33_ASAP7_75t_R register___U1013 ( .A(register__n202), .Y(register__n217) );
  INVxp33_ASAP7_75t_R register___U1014 ( .A(register__n202), .Y(register__n218) );
  INVxp33_ASAP7_75t_R register___U1015 ( .A(register__n203), .Y(register__n219) );
  INVxp33_ASAP7_75t_R register___U1016 ( .A(register__n203), .Y(register__n220) );
  INVxp33_ASAP7_75t_R register___U1017 ( .A(register__n203), .Y(register__n221) );
  AND2x2_ASAP7_75t_R register___U1018 ( .A(register__n12503), .B(register__n7684), .Y(register__n6302) );
  HB1xp67_ASAP7_75t_R register___U1019 ( .A(register__n218), .Y(register__n11819) );
  BUFx4f_ASAP7_75t_R register___U1020 ( .A(register__n3363), .Y(register__n3389) );
  INVxp67_ASAP7_75t_R register___U1021 ( .A(register__n11819), .Y(register__n1111) );
  INVxp67_ASAP7_75t_R register___U1022 ( .A(register__n11899), .Y(register__n11898) );
  CKINVDCx10_ASAP7_75t_R register___U1023 ( .A(register__n3734), .Y(register__n11896) );
  INVx6_ASAP7_75t_R register___U1024 ( .A(register__n11897), .Y(register__n3151) );
  BUFx2_ASAP7_75t_R register___U1025 ( .A(register__n6302), .Y(register__n11818) );
  BUFx3_ASAP7_75t_R register___U1026 ( .A(register__n6302), .Y(register__n3363) );
  INVx1_ASAP7_75t_R register___U1027 ( .A(write_data[27]), .Y(register__net63054) );
  BUFx4f_ASAP7_75t_R register___U1028 ( .A(register__n12224), .Y(register__n12206) );
  INVx2_ASAP7_75t_R register___U1029 ( .A(register__n12217), .Y(register__n12201) );
  BUFx2_ASAP7_75t_R register___U1030 ( .A(register__n5034), .Y(register__n12105) );
  INVx1_ASAP7_75t_R register___U1031 ( .A(register__n5034), .Y(register__n12083) );
  INVx1_ASAP7_75t_R register___U1032 ( .A(register__n12102), .Y(register__n12089) );
  INVx1_ASAP7_75t_R register___U1033 ( .A(register__n12106), .Y(register__n12092) );
  INVx1_ASAP7_75t_R register___U1034 ( .A(register__n12101), .Y(register__n12088) );
  INVx2_ASAP7_75t_R register___U1035 ( .A(register__n12105), .Y(register__n12091) );
  INVx2_ASAP7_75t_R register___U1036 ( .A(register__net88760), .Y(register__C6422_net60329) );
  OAI21x1_ASAP7_75t_R register___U1037 ( .A1(register__n2013), .A2(register__n2423), .B(register__n2448), .Y(register__n2443) );
  AND2x2_ASAP7_75t_R register___U1038 ( .A(register__n10838), .B(register__n7976), .Y(register__n1297) );
  NAND2x1_ASAP7_75t_R register___U1039 ( .A(register__n224), .B(register__n7300), .Y(register__n223) );
  AND4x1_ASAP7_75t_R register___U1040 ( .A(register__n1434), .B(register__n7929), .C(register__n7262), .D(register__n5588), .Y(
        n224) );
  HB1xp67_ASAP7_75t_R register___U1041 ( .A(register__n3741), .Y(register__n3740) );
  AOI22xp33_ASAP7_75t_R register___U1042 ( .A1(register__n1025), .A2(register__n1058), .B1(register__n1026), .B2(register__n1140), 
        .Y(register__n13173) );
  INVx5_ASAP7_75t_R register___U1043 ( .A(register__net63154), .Y(register__net140684) );
  INVx3_ASAP7_75t_R register___U1044 ( .A(register__net112808), .Y(register__net63154) );
  INVxp67_ASAP7_75t_R register___U1045 ( .A(write_data[25]), .Y(register__net112808) );
  AOI211xp5_ASAP7_75t_R register___U1046 ( .A1(register__n12521), .A2(register__n12517), .B(register__n747), .C(register__n746), 
        .Y(register__net61367) );
  NOR2x1_ASAP7_75t_R register___U1047 ( .A(register__n4964), .B(register__n4965), .Y(register__n747) );
  INVx1_ASAP7_75t_R register___U1048 ( .A(register__n13212), .Y(register__n225) );
  HB1xp67_ASAP7_75t_R register___U1049 ( .A(Reg_data[860]), .Y(register__n8211) );
  AND3x1_ASAP7_75t_R register___U1050 ( .A(register__n7638), .B(register__n7639), .C(register__n7640), .Y(register__n743) );
  AOI21xp5_ASAP7_75t_R register___U1051 ( .A1(register__C6423_net69526), .A2(register__net93508), .B(register__n2435), 
        .Y(register__n2455) );
  BUFx6f_ASAP7_75t_R register___U1052 ( .A(register__net144716), .Y(register__net146267) );
  HB1xp67_ASAP7_75t_R register___U1053 ( .A(register__n11147), .Y(register__n5024) );
  BUFx2_ASAP7_75t_R register___U1054 ( .A(register__n5024), .Y(register__n5023) );
  BUFx6f_ASAP7_75t_R register___U1055 ( .A(register__n3171), .Y(register__n3668) );
  BUFx6f_ASAP7_75t_R register___U1056 ( .A(register__n3187), .Y(register__n3171) );
  BUFx3_ASAP7_75t_R register___U1057 ( .A(register__n11982), .Y(register__n3187) );
  INVx2_ASAP7_75t_R register___U1058 ( .A(register__C6423_net61317), .Y(register__n1440) );
  AND2x2_ASAP7_75t_R register___U1059 ( .A(register__n389), .B(register__n11729), .Y(register__C6423_net61317) );
  INVxp67_ASAP7_75t_R register___U1060 ( .A(register__n1440), .Y(register__n1448) );
  INVxp67_ASAP7_75t_R register___U1061 ( .A(register__n1440), .Y(register__n1447) );
  INVxp67_ASAP7_75t_R register___U1062 ( .A(register__n1440), .Y(register__n1446) );
  INVxp67_ASAP7_75t_R register___U1063 ( .A(register__n1440), .Y(register__n1445) );
  INVxp33_ASAP7_75t_R register___U1064 ( .A(register__n1439), .Y(register__n1444) );
  BUFx6f_ASAP7_75t_R register___U1065 ( .A(register__n3340), .Y(register__n12391) );
  BUFx3_ASAP7_75t_R register___U1066 ( .A(register__n12392), .Y(register__n3340) );
  BUFx4f_ASAP7_75t_R register___U1067 ( .A(register__n2969), .Y(register__n2964) );
  BUFx4f_ASAP7_75t_R register___U1068 ( .A(register__net142724), .Y(register__net74013) );
  INVx1_ASAP7_75t_R register___U1069 ( .A(register__net142724), .Y(register__n1211) );
  INVx2_ASAP7_75t_R register___U1070 ( .A(register__n7114), .Y(register__n8578) );
  INVx3_ASAP7_75t_R register___U1071 ( .A(register__n3725), .Y(register__n12205) );
  INVx2_ASAP7_75t_R register___U1072 ( .A(register__n4025), .Y(register__n5927) );
  CKINVDCx20_ASAP7_75t_R register___U1073 ( .A(register__net98510), .Y(register__n227) );
  BUFx12_ASAP7_75t_R register___U1074 ( .A(register__net147145), .Y(register__net64390) );
  HB1xp67_ASAP7_75t_R register___U1075 ( .A(register__n13133), .Y(register__n3163) );
  AND2x6_ASAP7_75t_R register___U1076 ( .A(register__n11142), .B(register__n13), .Y(register__C6422_net60415) );
  BUFx2_ASAP7_75t_R register___U1077 ( .A(register__n2829), .Y(register__n11882) );
  AND2x4_ASAP7_75t_R register___U1078 ( .A(register__n10518), .B(register__n3407), .Y(register__n3908) );
  INVxp67_ASAP7_75t_R register___U1079 ( .A(register__n3025), .Y(register__n12370) );
  AND2x2_ASAP7_75t_R register___U1080 ( .A(register__n10518), .B(register__n12485), .Y(register__n1161) );
  INVx2_ASAP7_75t_R register___U1081 ( .A(register__n3264), .Y(register__n11861) );
  OAI22xp33_ASAP7_75t_R register___U1082 ( .A1(register__net64752), .A2(register__n2851), .B1(register__net89865), .B2(
        n3436), .Y(register__n228) );
  INVxp33_ASAP7_75t_R register___U1083 ( .A(register__n912), .Y(register__n229) );
  INVxp33_ASAP7_75t_R register___U1084 ( .A(register__n912), .Y(register__n230) );
  INVxp33_ASAP7_75t_R register___U1085 ( .A(register__n916), .Y(register__n930) );
  INVxp33_ASAP7_75t_R register___U1086 ( .A(register__n911), .Y(register__n920) );
  INVxp33_ASAP7_75t_R register___U1087 ( .A(register__n911), .Y(register__n919) );
  INVxp33_ASAP7_75t_R register___U1088 ( .A(register__n912), .Y(register__n921) );
  INVxp33_ASAP7_75t_R register___U1089 ( .A(register__n916), .Y(register__n929) );
  INVxp33_ASAP7_75t_R register___U1090 ( .A(register__n917), .Y(register__n931) );
  INVxp33_ASAP7_75t_R register___U1091 ( .A(register__n917), .Y(register__n932) );
  INVxp33_ASAP7_75t_R register___U1092 ( .A(register__n914), .Y(register__n926) );
  INVxp33_ASAP7_75t_R register___U1093 ( .A(register__n914), .Y(register__n925) );
  INVxp33_ASAP7_75t_R register___U1094 ( .A(register__n913), .Y(register__n923) );
  INVxp33_ASAP7_75t_R register___U1095 ( .A(register__n915), .Y(register__n928) );
  INVxp33_ASAP7_75t_R register___U1096 ( .A(register__n915), .Y(register__n927) );
  INVxp33_ASAP7_75t_R register___U1097 ( .A(register__net122579), .Y(register__n911) );
  INVxp33_ASAP7_75t_R register___U1098 ( .A(register__net122579), .Y(register__n917) );
  INVxp33_ASAP7_75t_R register___U1099 ( .A(register__net122579), .Y(register__n916) );
  INVxp67_ASAP7_75t_R register___U1100 ( .A(register__net122579), .Y(register__n912) );
  HB1xp67_ASAP7_75t_R register___U1101 ( .A(register__n8999), .Y(register__n8018) );
  HB1xp67_ASAP7_75t_R register___U1102 ( .A(register__n5082), .Y(register__n5081) );
  HB1xp67_ASAP7_75t_R register___U1103 ( .A(register__n3049), .Y(register__n3048) );
  BUFx4f_ASAP7_75t_R register___U1104 ( .A(register__net142380), .Y(register__net64360) );
  BUFx6f_ASAP7_75t_R register___U1105 ( .A(register__net117320), .Y(register__net64372) );
  NOR3x1_ASAP7_75t_R register___U1106 ( .A(register__n5333), .B(register__n9221), .C(register__n9219), .Y(register__n231) );
  BUFx6f_ASAP7_75t_R register___U1107 ( .A(register__n12388), .Y(register__n3025) );
  HB1xp67_ASAP7_75t_R register___U1108 ( .A(register__n12617), .Y(register__n4885) );
  HB1xp67_ASAP7_75t_R register___U1109 ( .A(register__net62718), .Y(register__net62716) );
  HB1xp67_ASAP7_75t_R register___U1110 ( .A(RegWrite), .Y(register__n1511) );
  INVx1_ASAP7_75t_R register___U1111 ( .A(register__n13104), .Y(register__n232) );
  AOI22xp33_ASAP7_75t_R register___U1112 ( .A1(register__n12044), .A2(register__n82), .B1(register__n664), .B2(register__n2799), 
        .Y(register__n12828) );
  NOR2xp67_ASAP7_75t_R register___U1113 ( .A(register__n11930), .B(register__n1069), .Y(register__n8601) );
  INVx1_ASAP7_75t_R register___U1114 ( .A(register__net122862), .Y(register__n_cell_124679_net155985) );
  HB1xp67_ASAP7_75t_R register___U1115 ( .A(register__n3117), .Y(register__n3116) );
  HB1xp67_ASAP7_75t_R register___U1116 ( .A(register__n11514), .Y(register__n4121) );
  AND2x2_ASAP7_75t_R register___U1117 ( .A(register__n1370), .B(register__n528), .Y(register__n9176) );
  INVx1_ASAP7_75t_R register___U1118 ( .A(register__n1440), .Y(register__n1449) );
  INVx3_ASAP7_75t_R register___U1119 ( .A(register__n4815), .Y(register__n12293) );
  BUFx3_ASAP7_75t_R register___U1120 ( .A(register__n12224), .Y(register__n3667) );
  INVx1_ASAP7_75t_R register___U1121 ( .A(register__n12950), .Y(register__n234) );
  HB1xp67_ASAP7_75t_R register___U1122 ( .A(register__n11597), .Y(register__n4471) );
  BUFx3_ASAP7_75t_R register___U1123 ( .A(register__net113802), .Y(register__net138040) );
  BUFx2_ASAP7_75t_R register___U1124 ( .A(register__n12494), .Y(register__n11762) );
  AOI22xp33_ASAP7_75t_R register___U1125 ( .A1(register__net64374), .A2(register__n5721), .B1(register__n236), .B2(
        n1411), .Y(register__n12998) );
  CKINVDCx20_ASAP7_75t_R register___U1126 ( .A(register__net90657), .Y(register__n236) );
  NAND4xp75_ASAP7_75t_R register___U1127 ( .A(register__n8558), .B(register__n8557), .C(register__n6830), .D(register__n8559), 
        .Y(register__n237) );
  AO22x1_ASAP7_75t_R register___U1128 ( .A1(register__n9905), .A2(register__net91683), .B1(register__n6384), .B2(register__n1358), 
        .Y(register__n10793) );
  AO22x1_ASAP7_75t_R register___U1129 ( .A1(register__n9660), .A2(register__n1867), .B1(register__net96692), .B2(register__n9989), 
        .Y(register__n10941) );
  AO22x1_ASAP7_75t_R register___U1130 ( .A1(register__net114112), .A2(register__n1867), .B1(register__net89401), .B2(
        net96692), .Y(register__n10809) );
  INVx2_ASAP7_75t_R register___U1131 ( .A(register__C6423_net60460), .Y(register__n709) );
  INVxp67_ASAP7_75t_R register___U1132 ( .A(register__n2874), .Y(register__n3912) );
  INVx1_ASAP7_75t_R register___U1133 ( .A(register__n3710), .Y(register__n984) );
  INVx1_ASAP7_75t_R register___U1134 ( .A(register__n12800), .Y(register__n238) );
  INVxp33_ASAP7_75t_R register___U1135 ( .A(register__net150876), .Y(register__n239) );
  AOI22x1_ASAP7_75t_R register___U1136 ( .A1(register__n12221), .A2(register__net130482), .B1(register__n397), .B2(
        net73055), .Y(register__n12647) );
  AO22x1_ASAP7_75t_R register___U1137 ( .A1(register__net62704), .A2(register__n346), .B1(register__n241), .B2(register__n337), 
        .Y(register__n240) );
  CKINVDCx20_ASAP7_75t_R register___U1138 ( .A(register__n8779), .Y(register__n241) );
  INVx1_ASAP7_75t_R register___U1139 ( .A(register__n336), .Y(register__n346) );
  NOR2xp67_ASAP7_75t_R register___U1140 ( .A(register__n7580), .B(register__n817), .Y(register__n621) );
  HB1xp67_ASAP7_75t_R register___U1141 ( .A(register__n10526), .Y(register__n5128) );
  INVx1_ASAP7_75t_R register___U1142 ( .A(register__n2838), .Y(register__n3752) );
  INVx1_ASAP7_75t_R register___U1143 ( .A(register__n1345), .Y(register__n1351) );
  HB1xp67_ASAP7_75t_R register___U1144 ( .A(register__n4219), .Y(register__n4218) );
  NAND2xp33_ASAP7_75t_R register___U1145 ( .A(register__n1851), .B(register__n606), .Y(register__n243) );
  NAND2xp5_ASAP7_75t_R register___U1146 ( .A(register__n242), .B(register__n243), .Y(read_reg_data_1[22]) );
  INVxp33_ASAP7_75t_R register___U1147 ( .A(register__n12383), .Y(register__n606) );
  NOR2xp67_ASAP7_75t_R register___U1148 ( .A(register__n570), .B(register__n571), .Y(register__n761) );
  BUFx2_ASAP7_75t_R register___U1149 ( .A(register__n10517), .Y(register__n3317) );
  BUFx3_ASAP7_75t_R register___U1150 ( .A(register__n3344), .Y(register__n3185) );
  INVx2_ASAP7_75t_R register___U1151 ( .A(register__net143769), .Y(register__n2147) );
  BUFx2_ASAP7_75t_R register___U1152 ( .A(register__net143769), .Y(register__net142724) );
  NOR2xp33_ASAP7_75t_R register___U1153 ( .A(register__n488), .B(register__n2470), .Y(register__n2472) );
  BUFx4f_ASAP7_75t_R register___U1154 ( .A(register__C6423_net61335), .Y(register__n2086) );
  INVx1_ASAP7_75t_R register___U1155 ( .A(register__n11975), .Y(register__n1471) );
  INVx2_ASAP7_75t_R register___U1156 ( .A(register__n11975), .Y(register__n11959) );
  INVxp33_ASAP7_75t_R register___U1157 ( .A(register__n11873), .Y(register__n987) );
  BUFx6f_ASAP7_75t_R register___U1158 ( .A(register__net110414), .Y(register__C6423_net69526) );
  INVx1_ASAP7_75t_R register___U1159 ( .A(register__n3793), .Y(register__n2127) );
  INVx1_ASAP7_75t_R register___U1160 ( .A(register__n2136), .Y(register__n1767) );
  AO22x1_ASAP7_75t_R register___U1161 ( .A1(register__n9742), .A2(register__net91683), .B1(register__n6609), .B2(
        net96692), .Y(register__n10770) );
  NAND2x1_ASAP7_75t_R register___U1162 ( .A(register__n6426), .B(register__n1290), .Y(register__n1289) );
  NAND2xp67_ASAP7_75t_R register___U1163 ( .A(register__n752), .B(register__n751), .Y(read_reg_data_1[25]) );
  BUFx2_ASAP7_75t_R register___U1164 ( .A(register__n3755), .Y(register__n5227) );
  HB1xp67_ASAP7_75t_R register___U1165 ( .A(register__n12482), .Y(register__n3755) );
  BUFx2_ASAP7_75t_R register___U1166 ( .A(register__n12482), .Y(register__n12480) );
  BUFx10_ASAP7_75t_R register___U1167 ( .A(register__n3002), .Y(register__n2986) );
  INVxp67_ASAP7_75t_R register___U1168 ( .A(register__n11709), .Y(register__n1085) );
  BUFx3_ASAP7_75t_R register___U1169 ( .A(register__n12165), .Y(register__n3541) );
  INVx2_ASAP7_75t_R register___U1170 ( .A(register__n1979), .Y(register__n1981) );
  INVx4_ASAP7_75t_R register___U1171 ( .A(register__n7633), .Y(register__n1951) );
  INVx2_ASAP7_75t_R register___U1172 ( .A(register__n11281), .Y(register__n9232) );
  INVxp67_ASAP7_75t_R register___U1173 ( .A(register__n3271), .Y(register__n6443) );
  HB1xp67_ASAP7_75t_R register___U1174 ( .A(rs2[4]), .Y(register__n244) );
  BUFx6f_ASAP7_75t_R register___U1175 ( .A(register__n739), .Y(register__n389) );
  BUFx2_ASAP7_75t_R register___U1176 ( .A(register__C6423_net60466), .Y(register__net131638) );
  NOR3xp33_ASAP7_75t_R register___U1177 ( .A(register__n10667), .B(register__n10669), .C(register__n10668), .Y(register__n864) );
  HB1xp67_ASAP7_75t_R register___U1178 ( .A(register__n2908), .Y(register__n2907) );
  INVx3_ASAP7_75t_R register___U1179 ( .A(register__n129), .Y(register__n481) );
  INVx2_ASAP7_75t_R register___U1180 ( .A(register__n762), .Y(register__net109849) );
  BUFx4_ASAP7_75t_R register___U1181 ( .A(register__n3604), .Y(register__n3513) );
  HB1xp67_ASAP7_75t_R register___U1182 ( .A(register__n883), .Y(register__net122599) );
  OAI22xp5_ASAP7_75t_R register___U1183 ( .A1(register__n245), .A2(register__n2021), .B1(register__n10116), .B2(register__n3426), 
        .Y(register__n525) );
  INVx13_ASAP7_75t_R register___U1184 ( .A(register__n2021), .Y(register__n2020) );
  HB1xp67_ASAP7_75t_R register___U1185 ( .A(register__n4778), .Y(register__n4777) );
  INVx4_ASAP7_75t_R register___U1186 ( .A(register__n12008), .Y(register__n11991) );
  OAI22xp33_ASAP7_75t_R register___U1187 ( .A1(register__net64008), .A2(register__n1973), .B1(register__net89397), .B2(
        n3408), .Y(register__n246) );
  NOR2xp67_ASAP7_75t_R register___U1188 ( .A(register__n1986), .B(register__n5389), .Y(register__n2747) );
  INVx1_ASAP7_75t_R register___U1189 ( .A(register__n1912), .Y(register__n1913) );
  AND2x2_ASAP7_75t_R register___U1190 ( .A(register__net109611), .B(register__n247), .Y(register__n414) );
  BUFx6f_ASAP7_75t_R register___U1191 ( .A(register__n3541), .Y(register__n3604) );
  INVxp33_ASAP7_75t_R register___U1192 ( .A(register__n260), .Y(register__n841) );
  INVxp67_ASAP7_75t_R register___U1193 ( .A(register__n5703), .Y(register__n2244) );
  NOR2xp33_ASAP7_75t_R register___U1194 ( .A(register__n11598), .B(register__n1274), .Y(register__n5703) );
  INVxp33_ASAP7_75t_R register___U1195 ( .A(register__net126578), .Y(register__net150873) );
  BUFx4f_ASAP7_75t_R register___U1196 ( .A(register__n11798), .Y(register__n11796) );
  NOR3xp33_ASAP7_75t_R register___U1197 ( .A(register__n248), .B(register__n249), .C(register__n250), .Y(register__n778) );
  NAND4xp75_ASAP7_75t_R register___U1198 ( .A(register__n6450), .B(register__n3835), .C(register__n6452), .D(register__n6451), 
        .Y(register__n248) );
  NAND4xp75_ASAP7_75t_R register___U1199 ( .A(register__n7910), .B(register__n7912), .C(register__n7911), .D(register__n7266), 
        .Y(register__n249) );
  NAND4xp25_ASAP7_75t_R register___U1200 ( .A(register__n3984), .B(register__n6147), .C(register__n8036), .D(register__n6149), 
        .Y(register__n250) );
  BUFx6f_ASAP7_75t_R register___U1201 ( .A(register__n2859), .Y(register__n3408) );
  INVx2_ASAP7_75t_R register___U1202 ( .A(register__n4120), .Y(register__n5233) );
  INVx6_ASAP7_75t_R register___U1203 ( .A(register__n6268), .Y(register__n12435) );
  INVx1_ASAP7_75t_R register___U1204 ( .A(register__n13130), .Y(register__n251) );
  INVx3_ASAP7_75t_R register___U1205 ( .A(register__n153), .Y(register__n482) );
  NOR2xp67_ASAP7_75t_R register___U1206 ( .A(register__n10641), .B(register__n2002), .Y(register__n252) );
  NOR2xp33_ASAP7_75t_R register___U1207 ( .A(register__n6212), .B(register__net112580), .Y(register__n254) );
  INVx2_ASAP7_75t_R register___U1208 ( .A(register__n9513), .Y(register__n10641) );
  HB1xp67_ASAP7_75t_R register___U1209 ( .A(register__n10642), .Y(register__n6212) );
  NOR2xp67_ASAP7_75t_R register___U1210 ( .A(register__n509), .B(register__n10), .Y(register__n2769) );
  AO22x1_ASAP7_75t_R register___U1211 ( .A1(register__n8527), .A2(register__n1867), .B1(register__n9433), .B2(register__n1351), 
        .Y(register__n10746) );
  AO22x1_ASAP7_75t_R register___U1212 ( .A1(register__n8765), .A2(register__n1867), .B1(register__n9987), .B2(register__net96692), 
        .Y(register__n10964) );
  HB1xp67_ASAP7_75t_R register___U1213 ( .A(register__n3027), .Y(register__n3026) );
  INVxp67_ASAP7_75t_R register___U1214 ( .A(register__n12993), .Y(register__n255) );
  AOI22xp33_ASAP7_75t_R register___U1215 ( .A1(register__n12242), .A2(register__n5721), .B1(register__n480), .B2(register__n1411), 
        .Y(register__n12993) );
  INVx1_ASAP7_75t_R register___U1216 ( .A(register__n2017), .Y(register__n1912) );
  BUFx6f_ASAP7_75t_R register___U1217 ( .A(register__n3667), .Y(register__n5442) );
  BUFx3_ASAP7_75t_R register___U1218 ( .A(register__n12223), .Y(register__n12222) );
  HB1xp67_ASAP7_75t_R register___U1219 ( .A(register__n12892), .Y(register__n3049) );
  HB1xp67_ASAP7_75t_R register___U1220 ( .A(register__n12897), .Y(register__n2908) );
  INVx2_ASAP7_75t_R register___U1221 ( .A(register__n5114), .Y(register__n7877) );
  NAND2xp33_ASAP7_75t_R register___U1222 ( .A(register__n8492), .B(register__net88727), .Y(register__n257) );
  NAND2xp33_ASAP7_75t_R register___U1223 ( .A(register__n256), .B(register__n257), .Y(register__n10797) );
  HB1xp67_ASAP7_75t_R register___U1224 ( .A(register__n10221), .Y(register__n8492) );
  HB1xp67_ASAP7_75t_R register___U1225 ( .A(register__n10797), .Y(register__n4810) );
  INVx1_ASAP7_75t_R register___U1226 ( .A(register__n5457), .Y(register__n258) );
  INVxp67_ASAP7_75t_R register___U1227 ( .A(register__n6497), .Y(register__n7949) );
  INVx1_ASAP7_75t_R register___U1228 ( .A(register__n11143), .Y(register__n1954) );
  OAI22xp5_ASAP7_75t_R register___U1229 ( .A1(register__net66316), .A2(register__n8585), .B1(register__n5350), .B2(
        n1687), .Y(read_reg_data_2[26]) );
  HB1xp67_ASAP7_75t_R register___U1230 ( .A(register__n11365), .Y(register__n8225) );
  HB1xp67_ASAP7_75t_R register___U1231 ( .A(register__n12618), .Y(register__n4006) );
  HB1xp67_ASAP7_75t_R register___U1232 ( .A(register__C6423_net61317), .Y(register__C6423_net72545) );
  AO22x1_ASAP7_75t_R register___U1233 ( .A1(register__n9603), .A2(register__C6423_net61318), .B1(register__n9427), .B2(
        C6423_net61317), .Y(register__n11230) );
  INVxp67_ASAP7_75t_R register___U1234 ( .A(register__C6423_net61317), .Y(register__n1439) );
  AND3x2_ASAP7_75t_R register___U1235 ( .A(register__n729), .B(IF_ID_rs1[2]), .C(register__n11143), .Y(
        n1012) );
  BUFx6f_ASAP7_75t_R register___U1236 ( .A(register__n12494), .Y(register__n3476) );
  NOR3xp33_ASAP7_75t_R register___U1237 ( .A(register__n6032), .B(register__n5116), .C(register__n8326), .Y(register__n259) );
  NAND2xp5_ASAP7_75t_R register___U1238 ( .A(register__n2189), .B(register__n2188), .Y(read_reg_data_2[27])
         );
  NAND2x2_ASAP7_75t_R register___U1239 ( .A(register__n655), .B(register__n818), .Y(register__n260) );
  INVx3_ASAP7_75t_R register___U1240 ( .A(register__net118635), .Y(register__n2342) );
  BUFx12f_ASAP7_75t_R register___U1241 ( .A(register__C6422_net70498), .Y(register__net118635) );
  OAI21xp33_ASAP7_75t_R register___U1242 ( .A1(register__n2345), .A2(register__n1420), .B(register__n2367), .Y(register__n2368)
         );
  OAI22xp33_ASAP7_75t_R register___U1243 ( .A1(register__n11932), .A2(register__n188), .B1(register__n9619), .B2(register__n217), 
        .Y(register__n261) );
  INVxp67_ASAP7_75t_R register___U1244 ( .A(register__n2015), .Y(register__n407) );
  INVxp67_ASAP7_75t_R register___U1245 ( .A(register__net150876), .Y(register__net150884) );
  HB1xp67_ASAP7_75t_R register___U1246 ( .A(register__n2875), .Y(register__n2874) );
  OAI22xp5_ASAP7_75t_R register___U1247 ( .A1(register__n1384), .A2(register__C6423_net72243), .B1(register__n1385), 
        .B2(register__n_cell_124679_net155985), .Y(register__n11397) );
  BUFx3_ASAP7_75t_R register___U1248 ( .A(register__net64398), .Y(register__net147145) );
  NAND3xp33_ASAP7_75t_R register___U1249 ( .A(register__n263), .B(register__n7018), .C(register__n7017), .Y(register__n1262) );
  NOR3xp33_ASAP7_75t_R register___U1250 ( .A(register__n1261), .B(register__n1262), .C(register__n1260), .Y(register__n2766) );
  NOR2x1_ASAP7_75t_R register___U1251 ( .A(register__n4822), .B(register__n11139), .Y(register__n1850) );
  BUFx2_ASAP7_75t_R register___U1252 ( .A(register__n11137), .Y(register__n4822) );
  AND2x2_ASAP7_75t_R register___U1253 ( .A(register__n1246), .B(register__n1323), .Y(register__n265) );
  AND3x1_ASAP7_75t_R register___U1254 ( .A(register__n265), .B(register__n4847), .C(register__n3209), .Y(register__n11260) );
  INVx3_ASAP7_75t_R register___U1255 ( .A(register__n5441), .Y(register__n11714) );
  HB1xp67_ASAP7_75t_R register___U1256 ( .A(register__n8230), .Y(register__n3209) );
  AO22x1_ASAP7_75t_R register___U1257 ( .A1(register__n9630), .A2(register__C6423_net69526), .B1(register__n10093), 
        .B2(register__net117890), .Y(register__n11236) );
  BUFx2_ASAP7_75t_R register___U1258 ( .A(register__n1951), .Y(register__n3711) );
  HB1xp67_ASAP7_75t_R register___U1259 ( .A(register__n11694), .Y(register__n5746) );
  INVx2_ASAP7_75t_R register___U1260 ( .A(write_data[13]), .Y(register__n12165) );
  INVx1_ASAP7_75t_R register___U1261 ( .A(register__n2086), .Y(register__n1903) );
  HB1xp67_ASAP7_75t_R register___U1262 ( .A(register__n11619), .Y(register__n5826) );
  OAI22xp33_ASAP7_75t_R register___U1263 ( .A1(register__n53), .A2(register__n7022), .B1(register__net61369), .B2(
        net64444), .Y(read_reg_data_1[10]) );
  HB1xp67_ASAP7_75t_R register___U1264 ( .A(register__n12766), .Y(register__n3780) );
  NOR2xp33_ASAP7_75t_R register___U1265 ( .A(register__n1687), .B(register__net64444), .Y(register__n2500) );
  HB1xp67_ASAP7_75t_R register___U1266 ( .A(register__n4243), .Y(register__n4242) );
  NOR2x1p5_ASAP7_75t_R register___U1267 ( .A(register__C6422_net59730), .B(register__net130666), .Y(register__n2372) );
  OAI22xp33_ASAP7_75t_R register___U1268 ( .A1(register__net66304), .A2(register__n6161), .B1(register__n12065), .B2(
        n1687), .Y(read_reg_data_2[8]) );
  HB1xp67_ASAP7_75t_R register___U1269 ( .A(register__n3272), .Y(register__n3271) );
  AND2x6_ASAP7_75t_R register___U1270 ( .A(register__n877), .B(register__n820), .Y(register__C6423_net61340) );
  INVx1_ASAP7_75t_R register___U1271 ( .A(register__n11050), .Y(register__n7304) );
  INVx2_ASAP7_75t_R register___U1272 ( .A(register__n11755), .Y(register__n1006) );
  NAND2x2_ASAP7_75t_R register___U1273 ( .A(register__n12483), .B(register__n1118), .Y(register__n2167) );
  INVxp67_ASAP7_75t_R register___U1274 ( .A(register__n3492), .Y(register__n8684) );
  HB1xp67_ASAP7_75t_R register___U1275 ( .A(register__n3493), .Y(register__n3492) );
  BUFx3_ASAP7_75t_R register___U1276 ( .A(register__net123880), .Y(register__net123879) );
  CKINVDCx6p67_ASAP7_75t_R register___U1277 ( .A(register__C6423_net60458), .Y(register__net130175) );
  INVx4_ASAP7_75t_R register___U1278 ( .A(register__n3171), .Y(register__n11954) );
  BUFx4f_ASAP7_75t_R register___U1279 ( .A(register__n11971), .Y(register__n3457) );
  INVx2_ASAP7_75t_R register___U1280 ( .A(register__n11954), .Y(register__n7611) );
  INVx2_ASAP7_75t_R register___U1281 ( .A(register__n3457), .Y(register__n11956) );
  HB1xp67_ASAP7_75t_R register___U1282 ( .A(register__n12673), .Y(register__n4420) );
  OAI22xp33_ASAP7_75t_R register___U1283 ( .A1(register__n11958), .A2(register__n109), .B1(register__n8787), .B2(register__n3451), 
        .Y(register__n266) );
  INVx1_ASAP7_75t_R register___U1284 ( .A(register__n10714), .Y(register__n267) );
  INVx5_ASAP7_75t_R register___U1285 ( .A(register__C6423_net60462), .Y(register__n2014) );
  HB1xp67_ASAP7_75t_R register___U1286 ( .A(register__n11465), .Y(register__n5600) );
  HB1xp67_ASAP7_75t_R register___U1287 ( .A(register__n13120), .Y(register__n3294) );
  BUFx6f_ASAP7_75t_R register___U1288 ( .A(register__n11780), .Y(register__n3302) );
  BUFx6f_ASAP7_75t_R register___U1289 ( .A(register__n3732), .Y(register__n12237) );
  OAI22xp5_ASAP7_75t_R register___U1290 ( .A1(register__n2123), .A2(register__net150044), .B1(register__n2124), .B2(
        n2023), .Y(register__n11401) );
  BUFx4f_ASAP7_75t_R register___U1291 ( .A(register__net117657), .Y(register__net88572) );
  INVx1_ASAP7_75t_R register___U1292 ( .A(register__n359), .Y(register__n360) );
  INVx6_ASAP7_75t_R register___U1293 ( .A(register__n2014), .Y(register__n2015) );
  BUFx2_ASAP7_75t_R register___U1294 ( .A(register__n7306), .Y(register__n4609) );
  INVxp67_ASAP7_75t_R register___U1295 ( .A(register__n4607), .Y(register__n7306) );
  BUFx3_ASAP7_75t_R register___U1296 ( .A(register__n11798), .Y(register__n11790) );
  OAI21xp33_ASAP7_75t_R register___U1297 ( .A1(register__n2332), .A2(register__n260), .B(register__n15), .Y(register__n2356) );
  BUFx3_ASAP7_75t_R register___U1298 ( .A(register__net64864), .Y(register__net143364) );
  INVx5_ASAP7_75t_R register___U1299 ( .A(write_data[5]), .Y(register__net64864) );
  BUFx4f_ASAP7_75t_R register___U1300 ( .A(register__net143364), .Y(register__net64884) );
  AND2x2_ASAP7_75t_R register___U1301 ( .A(register__n7020), .B(register__n11729), .Y(register__n268) );
  NAND2xp67_ASAP7_75t_R register___U1302 ( .A(register__n9365), .B(register__n840), .Y(register__n1515) );
  NAND2xp5_ASAP7_75t_R register___U1303 ( .A(register__n840), .B(register__net89777), .Y(register__n2401) );
  INVxp33_ASAP7_75t_R register___U1304 ( .A(register__n2010), .Y(register__n2011) );
  NOR3x1_ASAP7_75t_R register___U1305 ( .A(register__n6027), .B(register__n9207), .C(register__n9206), .Y(register__n269) );
  BUFx3_ASAP7_75t_R register___U1306 ( .A(register__n883), .Y(register__net113802) );
  BUFx2_ASAP7_75t_R register___U1307 ( .A(register__n2999), .Y(register__n2998) );
  INVx1_ASAP7_75t_R register___U1308 ( .A(register__n13086), .Y(register__n270) );
  NOR3xp33_ASAP7_75t_R register___U1309 ( .A(register__n10812), .B(register__n4164), .C(register__n10811), .Y(register__n271) );
  NOR2x1_ASAP7_75t_R register___U1310 ( .A(register__n8639), .B(register__n272), .Y(register__n10801) );
  INVxp67_ASAP7_75t_R register___U1311 ( .A(register__n271), .Y(register__n272) );
  BUFx2_ASAP7_75t_R register___U1312 ( .A(register__n10813), .Y(register__n4164) );
  INVx1_ASAP7_75t_R register___U1313 ( .A(register__n11154), .Y(register__n1760) );
  AOI22xp33_ASAP7_75t_R register___U1314 ( .A1(register__n3347), .A2(register__n5721), .B1(register__n553), .B2(register__n1411), 
        .Y(register__n12989) );
  BUFx12f_ASAP7_75t_R register___U1315 ( .A(register__n5349), .Y(register__n4198) );
  INVx1_ASAP7_75t_R register___U1316 ( .A(register__n3177), .Y(register__n2274) );
  HB1xp67_ASAP7_75t_R register___U1317 ( .A(register__n12224), .Y(register__n12223) );
  INVx1_ASAP7_75t_R register___U1318 ( .A(register__n13078), .Y(register__n273) );
  HB1xp67_ASAP7_75t_R register___U1319 ( .A(register__n13122), .Y(register__n2875) );
  HB1xp67_ASAP7_75t_R register___U1320 ( .A(Reg_data[13]), .Y(register__n8999) );
  INVx2_ASAP7_75t_R register___U1321 ( .A(register__n9523), .Y(register__n10760) );
  INVx5_ASAP7_75t_R register___U1322 ( .A(register__net113802), .Y(register__C6423_net72243) );
  AOI22xp33_ASAP7_75t_R register___U1323 ( .A1(register__n12331), .A2(register__n11783), .B1(register__n274), .B2(register__n1767), .Y(register__n12899) );
  CKINVDCx20_ASAP7_75t_R register___U1324 ( .A(register__n9971), .Y(register__n274) );
  INVx3_ASAP7_75t_R register___U1325 ( .A(register__n12331), .Y(register__n12318) );
  HB1xp67_ASAP7_75t_R register___U1326 ( .A(register__n2843), .Y(register__n11783) );
  AND2x4_ASAP7_75t_R register___U1327 ( .A(register__n11719), .B(register__n7020), .Y(register__C6423_net61326) );
  AND2x6_ASAP7_75t_R register___U1328 ( .A(register__n11149), .B(register__n11151), .Y(register__net126625) );
  CKINVDCx6p67_ASAP7_75t_R register___U1329 ( .A(register__n275), .Y(register__net93569) );
  INVxp67_ASAP7_75t_R register___U1330 ( .A(register__n1106), .Y(register__n308) );
  INVx1_ASAP7_75t_R register___U1331 ( .A(register__n308), .Y(register__n309) );
  CKINVDCx8_ASAP7_75t_R register___U1332 ( .A(register__C6423_net61325), .Y(register__n277) );
  INVxp67_ASAP7_75t_R register___U1333 ( .A(register__n13178), .Y(register__n6997) );
  INVxp67_ASAP7_75t_R register___U1334 ( .A(register__n12491), .Y(register__n3500) );
  INVx2_ASAP7_75t_R register___U1335 ( .A(register__n2849), .Y(register__n3835) );
  INVx1_ASAP7_75t_R register___U1336 ( .A(IF_ID_rs1[2]), .Y(register__n4490) );
  INVxp33_ASAP7_75t_R register___U1337 ( .A(register__n1239), .Y(register__n1240) );
  INVxp67_ASAP7_75t_R register___U1338 ( .A(register__net150876), .Y(register__net150896) );
  NAND4xp75_ASAP7_75t_R register___U1339 ( .A(register__n5698), .B(register__n5697), .C(register__n405), .D(register__n4328), .Y(
        n279) );
  NOR2xp33_ASAP7_75t_R register___U1340 ( .A(register__n2591), .B(register__n2615), .Y(register__n2617) );
  NOR2xp33_ASAP7_75t_R register___U1341 ( .A(register__n2622), .B(register__n545), .Y(register__n2623) );
  AND2x2_ASAP7_75t_R register___U1342 ( .A(register__n1224), .B(register__n1613), .Y(register__n280) );
  AND3x1_ASAP7_75t_R register___U1343 ( .A(register__n4337), .B(register__n280), .C(register__n5741), .Y(register__n11299) );
  INVxp67_ASAP7_75t_R register___U1344 ( .A(register__n9169), .Y(register__n5741) );
  AND4x2_ASAP7_75t_R register___U1345 ( .A(register__n7938), .B(register__n4185), .C(register__n7937), .D(register__n2224), .Y(
        n10974) );
  INVx2_ASAP7_75t_R register___U1346 ( .A(register__n3066), .Y(register__n7938) );
  HB1xp67_ASAP7_75t_R register___U1347 ( .A(register__n3300), .Y(register__n12379) );
  BUFx2_ASAP7_75t_R register___U1348 ( .A(register__n12392), .Y(register__n3342) );
  INVx1_ASAP7_75t_R register___U1349 ( .A(register__n13181), .Y(register__n282) );
  BUFx2_ASAP7_75t_R register___U1350 ( .A(register__net136186), .Y(register__net63028) );
  INVx1_ASAP7_75t_R register___U1351 ( .A(register__n12928), .Y(register__n283) );
  BUFx2_ASAP7_75t_R register___U1352 ( .A(register__C6423_net68950), .Y(register__C6423_net68948) );
  NOR3xp33_ASAP7_75t_R register___U1353 ( .A(register__n4027), .B(register__n4029), .C(register__n3920), .Y(register__n2797) );
  HB1xp67_ASAP7_75t_R register___U1354 ( .A(register__n4030), .Y(register__n4029) );
  INVx3_ASAP7_75t_R register___U1355 ( .A(register__n127), .Y(register__n285) );
  NOR2xp67_ASAP7_75t_R register___U1356 ( .A(register__n11557), .B(register__n1165), .Y(register__n286) );
  AND2x2_ASAP7_75t_R register___U1357 ( .A(register__n4759), .B(register__n1757), .Y(register__n288) );
  AND3x1_ASAP7_75t_R register___U1358 ( .A(register__n288), .B(register__n794), .C(register__n7908), .Y(register__n11428) );
  AO22x1_ASAP7_75t_R register___U1359 ( .A1(register__n9889), .A2(register__net125170), .B1(register__n10313), .B2(register__n515), .Y(register__n11461) );
  OAI22xp33_ASAP7_75t_R register___U1360 ( .A1(register__n11963), .A2(register__n1961), .B1(register__n8795), .B2(register__n1533), .Y(register__n289) );
  HB1xp67_ASAP7_75t_R register___U1361 ( .A(register__n12495), .Y(register__n3793) );
  INVx3_ASAP7_75t_R register___U1362 ( .A(register__n11720), .Y(register__n2739) );
  BUFx2_ASAP7_75t_R register___U1363 ( .A(register__n6466), .Y(register__n290) );
  AND2x6_ASAP7_75t_R register___U1364 ( .A(register__n5048), .B(register__n11152), .Y(register__C6422_net60445) );
  INVxp67_ASAP7_75t_R register___U1365 ( .A(register__n11154), .Y(register__n5048) );
  INVx2_ASAP7_75t_R register___U1366 ( .A(register__n2909), .Y(register__n4272) );
  AND2x4_ASAP7_75t_R register___U1367 ( .A(register__n8337), .B(register__n11728), .Y(register__n1998) );
  OAI21xp5_ASAP7_75t_R register___U1368 ( .A1(register__net99656), .A2(register__n2648), .B(register__n2670), .Y(register__n2669)
         );
  NOR4xp75_ASAP7_75t_R register___U1369 ( .A(register__n4024), .B(register__n4023), .C(register__n10833), .D(register__n4022), 
        .Y(register__n10818) );
  BUFx3_ASAP7_75t_R register___U1370 ( .A(register__n10831), .Y(register__n4024) );
  BUFx3_ASAP7_75t_R register___U1371 ( .A(register__n10832), .Y(register__n4023) );
  HB1xp67_ASAP7_75t_R register___U1372 ( .A(register__n11001), .Y(register__n2999) );
  NOR4xp75_ASAP7_75t_R register___U1373 ( .A(register__n3935), .B(register__n3934), .C(register__n10607), .D(register__n10605), 
        .Y(register__n10589) );
  BUFx3_ASAP7_75t_R register___U1374 ( .A(register__n10606), .Y(register__n3934) );
  BUFx3_ASAP7_75t_R register___U1375 ( .A(register__n10608), .Y(register__n3935) );
  INVxp67_ASAP7_75t_R register___U1376 ( .A(register__n5611), .Y(register__n6699) );
  BUFx6f_ASAP7_75t_R register___U1377 ( .A(register__n3704), .Y(register__n3571) );
  INVx2_ASAP7_75t_R register___U1378 ( .A(register__net129787), .Y(register__n_cell_125074_net170535) );
  HB1xp67_ASAP7_75t_R register___U1379 ( .A(register__n12952), .Y(register__n3493) );
  BUFx12f_ASAP7_75t_R register___U1380 ( .A(register__net64478), .Y(register__net91939) );
  BUFx12f_ASAP7_75t_R register___U1381 ( .A(register__net120961), .Y(register__net138612) );
  BUFx12f_ASAP7_75t_R register___U1382 ( .A(register__n1999), .Y(register__net120961) );
  INVx1_ASAP7_75t_R register___U1383 ( .A(register__n13144), .Y(register__n291) );
  INVx1_ASAP7_75t_R register___U1384 ( .A(register__n11115), .Y(register__n292) );
  INVxp67_ASAP7_75t_R register___U1385 ( .A(register__n5318), .Y(register__n293) );
  INVxp33_ASAP7_75t_R register___U1386 ( .A(WB_rd[1]), .Y(register__n294) );
  INVx1_ASAP7_75t_R register___U1387 ( .A(register__n12835), .Y(register__n295) );
  INVx1_ASAP7_75t_R register___U1388 ( .A(WB_rd[1]), .Y(register__n9408) );
  AND2x4_ASAP7_75t_R register___U1389 ( .A(WB_rd[2]), .B(WB_rd[1]), .Y(
        n593) );
  BUFx3_ASAP7_75t_R register___U1390 ( .A(WB_rd[1]), .Y(register__n5301) );
  INVx1_ASAP7_75t_R register___U1391 ( .A(register__n12836), .Y(register__n296) );
  INVx1_ASAP7_75t_R register___U1392 ( .A(register__n12894), .Y(register__n297) );
  INVx2_ASAP7_75t_R register___U1393 ( .A(register__n3230), .Y(register__n7882) );
  INVxp33_ASAP7_75t_R register___U1394 ( .A(register__n260), .Y(register__n837) );
  INVxp33_ASAP7_75t_R register___U1395 ( .A(register__n260), .Y(register__n836) );
  INVxp67_ASAP7_75t_R register___U1396 ( .A(register__n4421), .Y(register__n7249) );
  NAND3x1_ASAP7_75t_R register___U1397 ( .A(register__n1177), .B(register__n8277), .C(register__n5618), .Y(register__n2280) );
  HB1xp67_ASAP7_75t_R register___U1398 ( .A(register__n12889), .Y(register__n7355) );
  HB1xp67_ASAP7_75t_R register___U1399 ( .A(register__n11559), .Y(register__n3031) );
  AOI222xp33_ASAP7_75t_R register___U1400 ( .A1(register__net109611), .A2(register__n9501), .B1(register__n1993), .B2(
        n8706), .C1(register__n831), .C2(register__n9473), .Y(register__n11157) );
  INVx2_ASAP7_75t_R register___U1401 ( .A(register__net109611), .Y(register__net127626) );
  INVx1_ASAP7_75t_R register___U1402 ( .A(register__n9501), .Y(register__n10532) );
  INVx1_ASAP7_75t_R register___U1403 ( .A(register__n9473), .Y(register__n10534) );
  HB1xp67_ASAP7_75t_R register___U1404 ( .A(register__n4602), .Y(register__n4601) );
  OAI22xp33_ASAP7_75t_R register___U1405 ( .A1(register__n12422), .A2(register__n1705), .B1(register__n10333), .B2(
        n1693), .Y(register__n298) );
  INVx1_ASAP7_75t_R register___U1406 ( .A(register__n13242), .Y(register__n299) );
  BUFx3_ASAP7_75t_R register___U1407 ( .A(register__net63054), .Y(register__net136186) );
  INVxp33_ASAP7_75t_R register___U1408 ( .A(register__n406), .Y(register__n300) );
  AO22x1_ASAP7_75t_R register___U1409 ( .A1(register__n3171), .A2(register__n4579), .B1(register__n301), .B2(register__n1120), 
        .Y(register__n384) );
  CKINVDCx20_ASAP7_75t_R register___U1410 ( .A(register__n9339), .Y(register__n301) );
  BUFx4f_ASAP7_75t_R register___U1411 ( .A(register__n6430), .Y(register__n3350) );
  BUFx4f_ASAP7_75t_R register___U1412 ( .A(register__n5498), .Y(register__n3937) );
  NAND2xp5_ASAP7_75t_R register___U1413 ( .A(register__n1551), .B(register__n1554), .Y(register__n910) );
  INVx2_ASAP7_75t_R register___U1414 ( .A(WB_rd[3]), .Y(register__n12502) );
  BUFx6f_ASAP7_75t_R register___U1415 ( .A(register__net121619), .Y(register__C6422_net70498) );
  AOI22xp33_ASAP7_75t_R register___U1416 ( .A1(register__n5198), .A2(register__net93569), .B1(register__n4181), .B2(
        C6423_net74857), .Y(register__n302) );
  HB1xp67_ASAP7_75t_R register___U1417 ( .A(register__n3541), .Y(register__n12162) );
  INVx2_ASAP7_75t_R register___U1418 ( .A(register__n4618), .Y(register__n8627) );
  AOI22x1_ASAP7_75t_R register___U1419 ( .A1(register__net64970), .A2(register__n303), .B1(register__n304), .B2(register__n305), 
        .Y(register__n12796) );
  CKINVDCx20_ASAP7_75t_R register___U1420 ( .A(register__n2220), .Y(register__n303) );
  CKINVDCx20_ASAP7_75t_R register___U1421 ( .A(register__n9937), .Y(register__n304) );
  CKINVDCx20_ASAP7_75t_R register___U1422 ( .A(register__n5685), .Y(register__n305) );
  CKINVDCx5p33_ASAP7_75t_R register___U1423 ( .A(register__net64970), .Y(register__net64936) );
  OAI22xp33_ASAP7_75t_R register___U1424 ( .A1(register__n12148), .A2(register__n895), .B1(register__n9742), .B2(register__n897), 
        .Y(register__n306) );
  INVx1_ASAP7_75t_R register___U1425 ( .A(register__n13129), .Y(register__n3872) );
  BUFx6f_ASAP7_75t_R register___U1426 ( .A(register__n12267), .Y(register__n12264) );
  HB1xp67_ASAP7_75t_R register___U1427 ( .A(register__n12915), .Y(register__n3027) );
  INVxp33_ASAP7_75t_R register___U1428 ( .A(register__n3022), .Y(register__n307) );
  BUFx5_ASAP7_75t_R register___U1429 ( .A(register__n475), .Y(register__n3022) );
  INVx1_ASAP7_75t_R register___U1430 ( .A(register__n12804), .Y(register__n310) );
  INVxp67_ASAP7_75t_R register___U1431 ( .A(register__n5976), .Y(register__n9165) );
  NOR2xp67_ASAP7_75t_R register___U1432 ( .A(register__n1575), .B(register__n425), .Y(register__n483) );
  INVx1_ASAP7_75t_R register___U1433 ( .A(register__net145304), .Y(register__n454) );
  OR3x1_ASAP7_75t_R register___U1434 ( .A(register__n3178), .B(register__n1309), .C(register__n3180), .Y(register__n311) );
  INVxp33_ASAP7_75t_R register___U1435 ( .A(register__n1441), .Y(register__n1450) );
  INVxp67_ASAP7_75t_R register___U1436 ( .A(register__n1441), .Y(register__n1452) );
  INVxp67_ASAP7_75t_R register___U1437 ( .A(register__n1441), .Y(register__n1451) );
  INVx2_ASAP7_75t_R register___U1438 ( .A(register__n5628), .Y(register__n9396) );
  INVx3_ASAP7_75t_R register___U1439 ( .A(register__net63046), .Y(register__net124970) );
  OAI22xp5_ASAP7_75t_R register___U1440 ( .A1(register__n53), .A2(register__n9180), .B1(register__net61369), .B2(register__n11942), .Y(read_reg_data_1[0]) );
  INVxp33_ASAP7_75t_R register___U1441 ( .A(register__n3071), .Y(register__n1589) );
  BUFx6f_ASAP7_75t_R register___U1442 ( .A(register__n5641), .Y(register__n11741) );
  OAI22xp33_ASAP7_75t_R register___U1443 ( .A1(register__net63012), .A2(register__n7327), .B1(register__n9842), .B2(
        n5044), .Y(register__n313) );
  AND2x2_ASAP7_75t_R register___U1444 ( .A(register__n389), .B(register__n7996), .Y(register__C6423_net60456) );
  INVx6_ASAP7_75t_R register___U1445 ( .A(register__C6423_net60456), .Y(register__net131654) );
  BUFx3_ASAP7_75t_R register___U1446 ( .A(register__net131654), .Y(register__C6423_net68482) );
  BUFx3_ASAP7_75t_R register___U1447 ( .A(register__net131654), .Y(register__n2013) );
  INVxp67_ASAP7_75t_R register___U1448 ( .A(register__n4546), .Y(register__n5375) );
  HB1xp67_ASAP7_75t_R register___U1449 ( .A(register__n12526), .Y(register__n4546) );
  INVx1_ASAP7_75t_R register___U1450 ( .A(register__n10517), .Y(register__n1747) );
  INVx1_ASAP7_75t_R register___U1451 ( .A(register__n10517), .Y(register__n1746) );
  BUFx2_ASAP7_75t_R register___U1452 ( .A(register__n861), .Y(register__net147583) );
  BUFx3_ASAP7_75t_R register___U1453 ( .A(register__n3158), .Y(register__n3157) );
  OAI22xp33_ASAP7_75t_R register___U1454 ( .A1(register__net63012), .A2(register__n3343), .B1(register__n9353), .B2(
        n3248), .Y(register__n314) );
  BUFx12f_ASAP7_75t_R register___U1455 ( .A(register__n12189), .Y(register__n3512) );
  BUFx6f_ASAP7_75t_R register___U1456 ( .A(register__n709), .Y(register__n714) );
  BUFx3_ASAP7_75t_R register___U1457 ( .A(register__n285), .Y(register__net147378) );
  INVxp67_ASAP7_75t_R register___U1458 ( .A(register__n4837), .Y(register__n12233) );
  HB1xp67_ASAP7_75t_R register___U1459 ( .A(register__net91920), .Y(register__net64968) );
  NOR2x1_ASAP7_75t_R register___U1460 ( .A(register__n1459), .B(register__n11496), .Y(register__n315) );
  NOR2x1_ASAP7_75t_R register___U1461 ( .A(register__n1458), .B(register__n316), .Y(register__n4178) );
  INVx2_ASAP7_75t_R register___U1462 ( .A(register__n315), .Y(register__n316) );
  NAND2xp5_ASAP7_75t_R register___U1463 ( .A(register__n2251), .B(register__n2797), .Y(register__n1459) );
  NAND3x1_ASAP7_75t_R register___U1464 ( .A(register__n8574), .B(register__n4230), .C(register__n8575), .Y(register__n317) );
  NAND2x1_ASAP7_75t_R register___U1465 ( .A(register__n2928), .B(register__n318), .Y(register__n1318) );
  INVx1_ASAP7_75t_R register___U1466 ( .A(register__n317), .Y(register__n318) );
  INVx2_ASAP7_75t_R register___U1467 ( .A(register__n4231), .Y(register__n8574) );
  INVx2_ASAP7_75t_R register___U1468 ( .A(register__n4233), .Y(register__n8575) );
  BUFx3_ASAP7_75t_R register___U1469 ( .A(register__n8573), .Y(register__n4230) );
  BUFx12f_ASAP7_75t_R register___U1470 ( .A(register__n2846), .Y(register__n11798) );
  INVx2_ASAP7_75t_R register___U1471 ( .A(register__n2950), .Y(register__n11817) );
  BUFx2_ASAP7_75t_R register___U1472 ( .A(register__net128430), .Y(register__net64984) );
  INVxp33_ASAP7_75t_R register___U1473 ( .A(register__n300), .Y(register__n410) );
  INVx2_ASAP7_75t_R register___U1474 ( .A(write_data[1]), .Y(register__n11982) );
  AOI22x1_ASAP7_75t_R register___U1475 ( .A1(register__n11966), .A2(register__n319), .B1(register__n320), .B2(register__n321), 
        .Y(register__n13387) );
  CKINVDCx20_ASAP7_75t_R register___U1476 ( .A(register__n11730), .Y(register__n319) );
  CKINVDCx20_ASAP7_75t_R register___U1477 ( .A(register__n10361), .Y(register__n320) );
  CKINVDCx20_ASAP7_75t_R register___U1478 ( .A(register__n1164), .Y(register__n321) );
  CKINVDCx5p33_ASAP7_75t_R register___U1479 ( .A(register__n11966), .Y(register__n11949) );
  AO22x1_ASAP7_75t_R register___U1480 ( .A1(register__net63042), .A2(register__n4270), .B1(register__n323), .B2(register__n11829), 
        .Y(register__n322) );
  CKINVDCx20_ASAP7_75t_R register___U1481 ( .A(register__n9840), .Y(register__n323) );
  AND2x6_ASAP7_75t_R register___U1482 ( .A(register__n11142), .B(register__n11151), .Y(register__net120912) );
  INVx1_ASAP7_75t_R register___U1483 ( .A(register__n12909), .Y(register__n324) );
  INVx1_ASAP7_75t_R register___U1484 ( .A(register__n12827), .Y(register__n325) );
  NAND2xp5_ASAP7_75t_R register___U1485 ( .A(register__n50), .B(register__n872), .Y(register__n530) );
  AO22x1_ASAP7_75t_R register___U1486 ( .A1(register__n6620), .A2(register__n77), .B1(register__n9935), .B2(register__n75), .Y(
        n10675) );
  AO22x1_ASAP7_75t_R register___U1487 ( .A1(register__n6897), .A2(register__n77), .B1(register__n9929), .B2(register__n75), .Y(
        n10970) );
  AO22x1_ASAP7_75t_R register___U1488 ( .A1(register__n6956), .A2(register__n77), .B1(register__n10471), .B2(register__n75), .Y(
        n10903) );
  AO22x1_ASAP7_75t_R register___U1489 ( .A1(register__net107859), .A2(register__n77), .B1(register__net89001), .B2(register__n75), 
        .Y(register__n11094) );
  BUFx6f_ASAP7_75t_R register___U1490 ( .A(register__n11851), .Y(register__n3426) );
  HB1xp67_ASAP7_75t_R register___U1491 ( .A(register__n3426), .Y(register__n4952) );
  CKINVDCx8_ASAP7_75t_R register___U1492 ( .A(register__n3324), .Y(register__n1092) );
  INVxp67_ASAP7_75t_R register___U1493 ( .A(register__n6781), .Y(register__n7894) );
  INVxp67_ASAP7_75t_R register___U1494 ( .A(register__n4007), .Y(register__n4856) );
  INVxp67_ASAP7_75t_R register___U1495 ( .A(register__n5160), .Y(register__n8312) );
  BUFx6f_ASAP7_75t_R register___U1496 ( .A(register__net100543), .Y(register__net100540) );
  BUFx6f_ASAP7_75t_R register___U1497 ( .A(register__net100543), .Y(register__net100542) );
  BUFx6f_ASAP7_75t_R register___U1498 ( .A(register__net148003), .Y(register__net64472) );
  BUFx6f_ASAP7_75t_R register___U1499 ( .A(register__C6423_net61340), .Y(register__net141083) );
  INVxp33_ASAP7_75t_R register___U1500 ( .A(register__n1979), .Y(register__n1983) );
  INVxp33_ASAP7_75t_R register___U1501 ( .A(register__n1979), .Y(register__n1982) );
  INVxp33_ASAP7_75t_R register___U1502 ( .A(register__n1979), .Y(register__n1980) );
  INVxp67_ASAP7_75t_R register___U1503 ( .A(register__n1984), .Y(register__n1527) );
  INVx3_ASAP7_75t_R register___U1504 ( .A(register__n1984), .Y(register__n1979) );
  BUFx6f_ASAP7_75t_R register___U1505 ( .A(register__n12336), .Y(register__n12335) );
  BUFx6f_ASAP7_75t_R register___U1506 ( .A(register__n12050), .Y(register__n4865) );
  INVx1_ASAP7_75t_R register___U1507 ( .A(register__n1503), .Y(register__n6467) );
  HB1xp67_ASAP7_75t_R register___U1508 ( .A(register__n1773), .Y(register__n11803) );
  BUFx12f_ASAP7_75t_R register___U1509 ( .A(register__net62850), .Y(register__net141520) );
  HB1xp67_ASAP7_75t_R register___U1510 ( .A(register__n13360), .Y(register__n4012) );
  BUFx3_ASAP7_75t_R register___U1511 ( .A(register__net109849), .Y(register__net128109) );
  INVxp67_ASAP7_75t_R register___U1512 ( .A(register__n4331), .Y(register__n7643) );
  INVxp67_ASAP7_75t_R register___U1513 ( .A(register__n12605), .Y(register__n6731) );
  INVx4_ASAP7_75t_R register___U1514 ( .A(register__n4031), .Y(register__n12151) );
  BUFx6f_ASAP7_75t_R register___U1515 ( .A(register__n12162), .Y(register__n3219) );
  OAI22xp5_ASAP7_75t_R register___U1516 ( .A1(register__n12143), .A2(register__n11862), .B1(register__n10108), .B2(
        n3382), .Y(register__n1688) );
  INVx6_ASAP7_75t_R register___U1517 ( .A(register__n3946), .Y(register__n11862) );
  NAND2xp5_ASAP7_75t_R register___U1518 ( .A(register__n19), .B(register__n530), .Y(read_reg_data_1[17]) );
  AOI222xp33_ASAP7_75t_R register___U1519 ( .A1(register__net109611), .A2(register__n10373), .B1(register__net131638), 
        .B2(register__n8282), .C1(register__n831), .C2(register__n10378), .Y(register__n11388) );
  INVx2_ASAP7_75t_R register___U1520 ( .A(register__n10765), .Y(register__n9158) );
  BUFx6f_ASAP7_75t_R register___U1521 ( .A(register__net63390), .Y(register__net143520) );
  HB1xp67_ASAP7_75t_R register___U1522 ( .A(register__n7052), .Y(register__n328) );
  AND3x1_ASAP7_75t_R register___U1523 ( .A(register__n9168), .B(register__n7299), .C(register__n7298), .Y(register__n329) );
  AND2x2_ASAP7_75t_R register___U1524 ( .A(register__n4900), .B(register__n329), .Y(register__n11175) );
  BUFx6f_ASAP7_75t_R register___U1525 ( .A(register__n12206), .Y(register__n6404) );
  INVx4_ASAP7_75t_R register___U1526 ( .A(write_data[23]), .Y(register__net63390) );
  OAI22xp33_ASAP7_75t_R register___U1527 ( .A1(register__net62994), .A2(register__n1092), .B1(register__n6973), .B2(
        n3476), .Y(register__n330) );
  AND2x2_ASAP7_75t_R register___U1528 ( .A(register__n1429), .B(register__n6715), .Y(register__n331) );
  AND2x2_ASAP7_75t_R register___U1529 ( .A(register__n6714), .B(register__n331), .Y(register__n1259) );
  BUFx3_ASAP7_75t_R register___U1530 ( .A(register__n11993), .Y(register__n3593) );
  BUFx6f_ASAP7_75t_R register___U1531 ( .A(register__n12017), .Y(register__n11999) );
  CKINVDCx8_ASAP7_75t_R register___U1532 ( .A(register__C6423_net60466), .Y(register__n1995) );
  INVx3_ASAP7_75t_R register___U1533 ( .A(register__n3940), .Y(register__n3939) );
  NOR2x1p5_ASAP7_75t_R register___U1534 ( .A(register__n2127), .B(register__n3939), .Y(register__n12498) );
  HB1xp67_ASAP7_75t_R register___U1535 ( .A(register__n4422), .Y(register__n4421) );
  INVx2_ASAP7_75t_R register___U1536 ( .A(register__C6423_net60460), .Y(register__n710) );
  NAND2xp33_ASAP7_75t_R register___U1537 ( .A(register__n820), .B(register__n11729), .Y(register__n2157) );
  NAND2xp33_ASAP7_75t_R register___U1538 ( .A(register__n10205), .B(register__n285), .Y(register__n1378) );
  INVx2_ASAP7_75t_R register___U1539 ( .A(register__n4559), .Y(register__n6420) );
  INVxp67_ASAP7_75t_R register___U1540 ( .A(register__n5749), .Y(register__n7281) );
  HB1xp67_ASAP7_75t_R register___U1541 ( .A(register__n5750), .Y(register__n5749) );
  BUFx12f_ASAP7_75t_R register___U1542 ( .A(register__n4745), .Y(register__n3844) );
  BUFx6f_ASAP7_75t_R register___U1543 ( .A(register__n12309), .Y(register__n4745) );
  INVx2_ASAP7_75t_R register___U1544 ( .A(n3), .Y(register__n12278) );
  INVxp67_ASAP7_75t_R register___U1545 ( .A(register__n8364), .Y(register__n9403) );
  HB1xp67_ASAP7_75t_R register___U1546 ( .A(register__n8365), .Y(register__n8364) );
  BUFx6f_ASAP7_75t_R register___U1547 ( .A(register__n3651), .Y(register__n3349) );
  HB1xp67_ASAP7_75t_R register___U1548 ( .A(register__n10728), .Y(register__n4243) );
  BUFx6f_ASAP7_75t_R register___U1549 ( .A(register__n4967), .Y(register__n3601) );
  BUFx3_ASAP7_75t_R register___U1550 ( .A(register__n2960), .Y(register__n11801) );
  INVxp67_ASAP7_75t_R register___U1551 ( .A(register__n5773), .Y(register__n6737) );
  HB1xp67_ASAP7_75t_R register___U1552 ( .A(register__n5774), .Y(register__n5773) );
  AO22x1_ASAP7_75t_R register___U1553 ( .A1(register__net62876), .A2(register__n1603), .B1(register__n333), .B2(register__n2935), 
        .Y(register__n332) );
  CKINVDCx20_ASAP7_75t_R register___U1554 ( .A(register__net88756), .Y(register__n333) );
  INVx2_ASAP7_75t_R register___U1555 ( .A(register__net62876), .Y(register__net62840) );
  INVx1_ASAP7_75t_R register___U1556 ( .A(register__n3022), .Y(register__n1603) );
  CKINVDCx10_ASAP7_75t_R register___U1557 ( .A(register__C6422_net59544), .Y(register__n1691) );
  BUFx6f_ASAP7_75t_R register___U1558 ( .A(register__n3158), .Y(register__n3156) );
  BUFx6f_ASAP7_75t_R register___U1559 ( .A(register__n3187), .Y(register__n3158) );
  NAND2xp33_ASAP7_75t_R register___U1560 ( .A(register__n278), .B(register__n876), .Y(register__n1470) );
  INVxp33_ASAP7_75t_R register___U1561 ( .A(register__n875), .Y(register__n876) );
  BUFx6f_ASAP7_75t_R register___U1562 ( .A(register__n3260), .Y(register__n3259) );
  INVx1_ASAP7_75t_R register___U1563 ( .A(register__n102), .Y(register__n335) );
  INVx1_ASAP7_75t_R register___U1564 ( .A(register__n102), .Y(register__n338) );
  INVx4_ASAP7_75t_R register___U1565 ( .A(register__n337), .Y(register__n342) );
  INVx1_ASAP7_75t_R register___U1566 ( .A(register__n340), .Y(register__n343) );
  INVx1_ASAP7_75t_R register___U1567 ( .A(register__n341), .Y(register__n344) );
  INVx1_ASAP7_75t_R register___U1568 ( .A(register__n339), .Y(register__n345) );
  HB1xp67_ASAP7_75t_R register___U1569 ( .A(register__n3286), .Y(register__n3285) );
  AND2x6_ASAP7_75t_R register___U1570 ( .A(register__n448), .B(register__n312), .Y(register__net126316) );
  AO22x1_ASAP7_75t_R register___U1571 ( .A1(register__n9871), .A2(register__n1909), .B1(register__n10285), .B2(register__n1579), 
        .Y(register__n11033) );
  HB1xp67_ASAP7_75t_R register___U1572 ( .A(register__n13217), .Y(register__n5571) );
  HB1xp67_ASAP7_75t_R register___U1573 ( .A(register__n13187), .Y(register__n5768) );
  INVx6_ASAP7_75t_R register___U1574 ( .A(register__net63266), .Y(register__net103248) );
  INVx6_ASAP7_75t_R register___U1575 ( .A(register__net127751), .Y(register__net63266) );
  INVxp67_ASAP7_75t_R register___U1576 ( .A(register__n5013), .Y(register__n7086) );
  HB1xp67_ASAP7_75t_R register___U1577 ( .A(register__n5014), .Y(register__n5013) );
  INVxp67_ASAP7_75t_R register___U1578 ( .A(register__n4873), .Y(register__n6682) );
  HB1xp67_ASAP7_75t_R register___U1579 ( .A(register__n4874), .Y(register__n4873) );
  INVx1_ASAP7_75t_R register___U1580 ( .A(register__n4934), .Y(register__n8314) );
  INVxp33_ASAP7_75t_R register___U1581 ( .A(register__net64942), .Y(register__n1382) );
  INVx1_ASAP7_75t_R register___U1582 ( .A(register__net64942), .Y(register__net134980) );
  INVx6_ASAP7_75t_R register___U1583 ( .A(register__net127323), .Y(register__net64916) );
  BUFx6f_ASAP7_75t_R register___U1584 ( .A(register__net127323), .Y(register__net64960) );
  CKINVDCx6p67_ASAP7_75t_R register___U1585 ( .A(register__net64924), .Y(register__net127323) );
  CKINVDCx8_ASAP7_75t_R register___U1586 ( .A(register__net91921), .Y(register__net64924) );
  NAND2xp33_ASAP7_75t_R register___U1587 ( .A(register__n348), .B(register__n349), .Y(register__n10673) );
  NOR3xp33_ASAP7_75t_R register___U1588 ( .A(register__n31), .B(register__n4103), .C(register__n1373), .Y(register__n10656) );
  BUFx3_ASAP7_75t_R register___U1589 ( .A(register__n8784), .Y(register__n8783) );
  INVx1_ASAP7_75t_R register___U1590 ( .A(register__n4107), .Y(register__n1373) );
  AND2x2_ASAP7_75t_R register___U1591 ( .A(register__n154), .B(register__n5301), .Y(register__n9389) );
  XNOR2x2_ASAP7_75t_R register___U1592 ( .A(register__n1489), .B(register__n5301), .Y(register__n12519) );
  HB1xp67_ASAP7_75t_R register___U1593 ( .A(register__n6721), .Y(register__n5183) );
  INVx6_ASAP7_75t_R register___U1594 ( .A(register__n2829), .Y(register__n11881) );
  INVx1_ASAP7_75t_R register___U1595 ( .A(register__n11882), .Y(register__n1301) );
  OAI22xp5_ASAP7_75t_R register___U1596 ( .A1(register__net112762), .A2(register__n9155), .B1(register__net64966), .B2(
        n1687), .Y(read_reg_data_2[4]) );
  BUFx4f_ASAP7_75t_R register___U1597 ( .A(register__n5045), .Y(register__n4578) );
  BUFx6f_ASAP7_75t_R register___U1598 ( .A(register__C6423_net72238), .Y(register__net122601) );
  INVx1_ASAP7_75t_R register___U1599 ( .A(register__n10976), .Y(register__n350) );
  INVx1_ASAP7_75t_R register___U1600 ( .A(register__n12596), .Y(register__n351) );
  BUFx4f_ASAP7_75t_R register___U1601 ( .A(register__n3711), .Y(register__n3709) );
  INVx3_ASAP7_75t_R register___U1602 ( .A(register__n7674), .Y(register__n5124) );
  BUFx4f_ASAP7_75t_R register___U1603 ( .A(register__n3516), .Y(register__n3515) );
  INVx2_ASAP7_75t_R register___U1604 ( .A(register__n12362), .Y(register__n12347) );
  CKINVDCx8_ASAP7_75t_R register___U1605 ( .A(register__n5344), .Y(register__n12350) );
  BUFx2_ASAP7_75t_R register___U1606 ( .A(register__n12165), .Y(register__n12164) );
  OAI22xp33_ASAP7_75t_R register___U1607 ( .A1(register__net64422), .A2(register__n1092), .B1(register__net90401), .B2(
        n3918), .Y(register__n352) );
  HB1xp67_ASAP7_75t_R register___U1608 ( .A(register__n13297), .Y(register__n4887) );
  INVx2_ASAP7_75t_R register___U1609 ( .A(register__n2286), .Y(register__n11826) );
  BUFx4f_ASAP7_75t_R register___U1610 ( .A(register__n12050), .Y(register__n3837) );
  BUFx2_ASAP7_75t_R register___U1611 ( .A(register__n4865), .Y(register__n12034) );
  HB1xp67_ASAP7_75t_R register___U1612 ( .A(register__n13050), .Y(register__n5082) );
  HB1xp67_ASAP7_75t_R register___U1613 ( .A(register__net122862), .Y(register__net139882) );
  INVxp67_ASAP7_75t_R register___U1614 ( .A(register__n2884), .Y(register__n3440) );
  HB1xp67_ASAP7_75t_R register___U1615 ( .A(register__n2885), .Y(register__n2884) );
  HB1xp67_ASAP7_75t_R register___U1616 ( .A(register__n11636), .Y(register__n2885) );
  INVx4_ASAP7_75t_R register___U1617 ( .A(register__net138885), .Y(register__net63338) );
  NAND4xp75_ASAP7_75t_R register___U1618 ( .A(register__n7605), .B(register__n1421), .C(register__n7606), .D(register__n8578), 
        .Y(register__n509) );
  AO22x1_ASAP7_75t_R register___U1619 ( .A1(register__net63356), .A2(register__n4968), .B1(register__n355), .B2(register__n887), 
        .Y(register__n354) );
  CKINVDCx20_ASAP7_75t_R register___U1620 ( .A(register__n9415), .Y(register__n355) );
  INVx1_ASAP7_75t_R register___U1621 ( .A(register__n887), .Y(register__n901) );
  INVx1_ASAP7_75t_R register___U1622 ( .A(register__n12961), .Y(register__n356) );
  HB1xp67_ASAP7_75t_R register___U1623 ( .A(register__n11277), .Y(register__n3208) );
  INVx1_ASAP7_75t_R register___U1624 ( .A(register__n13069), .Y(register__n357) );
  BUFx6f_ASAP7_75t_R register___U1625 ( .A(register__net125365), .Y(register__C6423_net69198) );
  BUFx3_ASAP7_75t_R register___U1626 ( .A(register__n8235), .Y(register__n5255) );
  HB1xp67_ASAP7_75t_R register___U1627 ( .A(register__n10803), .Y(register__n5160) );
  INVx1_ASAP7_75t_R register___U1628 ( .A(register__n11056), .Y(register__n358) );
  HB1xp67_ASAP7_75t_R register___U1629 ( .A(register__n12666), .Y(register__n4422) );
  INVxp33_ASAP7_75t_R register___U1630 ( .A(register__net121558), .Y(register__net126578) );
  INVxp33_ASAP7_75t_R register___U1631 ( .A(register__n1998), .Y(register__net150878) );
  INVx3_ASAP7_75t_R register___U1632 ( .A(register__n1998), .Y(register__n2019) );
  BUFx12f_ASAP7_75t_R register___U1633 ( .A(register__n3451), .Y(register__n5504) );
  BUFx6f_ASAP7_75t_R register___U1634 ( .A(register__n1774), .Y(register__n3451) );
  NAND2xp67_ASAP7_75t_R register___U1635 ( .A(register__n10950), .B(register__n761), .Y(register__n359) );
  OAI22xp33_ASAP7_75t_R register___U1636 ( .A1(register__net64836), .A2(register__n1616), .B1(register__net90829), .B2(
        n3509), .Y(register__n361) );
  BUFx6f_ASAP7_75t_R register___U1637 ( .A(register__net142380), .Y(register__net142573) );
  BUFx6f_ASAP7_75t_R register___U1638 ( .A(register__net64398), .Y(register__net142380) );
  INVx1_ASAP7_75t_R register___U1639 ( .A(register__n653), .Y(register__n1953) );
  INVx1_ASAP7_75t_R register___U1640 ( .A(register__n653), .Y(register__n597) );
  INVxp33_ASAP7_75t_R register___U1641 ( .A(register__n1299), .Y(register__n726) );
  BUFx2_ASAP7_75t_R register___U1642 ( .A(register__n12191), .Y(register__n3375) );
  INVx2_ASAP7_75t_R register___U1643 ( .A(register__n4470), .Y(register__n5706) );
  INVx4_ASAP7_75t_R register___U1644 ( .A(register__n9521), .Y(register__n11060) );
  INVx6_ASAP7_75t_R register___U1645 ( .A(register__net143694), .Y(register__net63994) );
  INVxp33_ASAP7_75t_R register___U1646 ( .A(register__n4837), .Y(register__n3443) );
  BUFx2_ASAP7_75t_R register___U1647 ( .A(register__n2863), .Y(register__n2862) );
  HB1xp67_ASAP7_75t_R register___U1648 ( .A(register__n11318), .Y(register__n2863) );
  INVx1_ASAP7_75t_R register___U1649 ( .A(register__n13085), .Y(register__n362) );
  AO22x1_ASAP7_75t_R register___U1650 ( .A1(register__net148409), .A2(register__n1593), .B1(register__net113148), .B2(
        n1991), .Y(register__n363) );
  INVx1_ASAP7_75t_R register___U1651 ( .A(register__n2139), .Y(register__n1991) );
  INVx2_ASAP7_75t_R register___U1652 ( .A(register__n1991), .Y(register__n1593) );
  NOR2xp67_ASAP7_75t_R register___U1653 ( .A(register__n1997), .B(register__n11064), .Y(register__n786) );
  INVx4_ASAP7_75t_R register___U1654 ( .A(register__n10419), .Y(register__n11064) );
  INVxp67_ASAP7_75t_R register___U1655 ( .A(register__n5087), .Y(register__n6741) );
  HB1xp67_ASAP7_75t_R register___U1656 ( .A(register__n5088), .Y(register__n5087) );
  HB1xp67_ASAP7_75t_R register___U1657 ( .A(register__n12741), .Y(register__n3395) );
  AND2x2_ASAP7_75t_R register___U1658 ( .A(register__n820), .B(register__n1107), .Y(register__net122579) );
  INVx5_ASAP7_75t_R register___U1659 ( .A(register__n11726), .Y(register__n7020) );
  BUFx6f_ASAP7_75t_R register___U1660 ( .A(register__net141459), .Y(register__net64780) );
  BUFx12f_ASAP7_75t_R register___U1661 ( .A(register__net127692), .Y(register__net64790) );
  INVx3_ASAP7_75t_R register___U1662 ( .A(write_data[6]), .Y(register__net64818) );
  INVx2_ASAP7_75t_R register___U1663 ( .A(write_data[24]), .Y(register__n667) );
  INVx1_ASAP7_75t_R register___U1664 ( .A(register__n10930), .Y(register__n364) );
  INVx2_ASAP7_75t_R register___U1665 ( .A(register__n5607), .Y(register__n6697) );
  INVx1_ASAP7_75t_R register___U1666 ( .A(register__n13051), .Y(register__n365) );
  CKINVDCx8_ASAP7_75t_R register___U1667 ( .A(register__net143363), .Y(register__net64832) );
  BUFx12f_ASAP7_75t_R register___U1668 ( .A(register__net64864), .Y(register__net143363) );
  INVx6_ASAP7_75t_R register___U1669 ( .A(register__net64832), .Y(register__net102927) );
  BUFx4f_ASAP7_75t_R register___U1670 ( .A(register__n12351), .Y(register__n12360) );
  OAI21xp5_ASAP7_75t_R register___U1671 ( .A1(register__net99656), .A2(register__n2381), .B(register__n2401), .Y(register__n2400)
         );
  INVx6_ASAP7_75t_R register___U1672 ( .A(register__n12351), .Y(register__n12339) );
  NOR2xp67_ASAP7_75t_R register___U1673 ( .A(register__n24), .B(register__n2394), .Y(register__n2397) );
  INVx1_ASAP7_75t_R register___U1674 ( .A(register__n594), .Y(register__n1510) );
  BUFx3_ASAP7_75t_R register___U1675 ( .A(register__n3511), .Y(register__n3510) );
  HB1xp67_ASAP7_75t_R register___U1676 ( .A(register__n12030), .Y(register__n3665) );
  INVx1_ASAP7_75t_R register___U1677 ( .A(register__n10553), .Y(register__n7671) );
  INVxp67_ASAP7_75t_R register___U1678 ( .A(register__n2016), .Y(register__n2017) );
  BUFx12f_ASAP7_75t_R register___U1679 ( .A(register__net117658), .Y(register__net117657) );
  NOR2xp33_ASAP7_75t_R register___U1680 ( .A(register__n1987), .B(register__n10915), .Y(register__n2752) );
  BUFx3_ASAP7_75t_R register___U1681 ( .A(register__n7686), .Y(register__n4964) );
  BUFx6f_ASAP7_75t_R register___U1682 ( .A(register__n11883), .Y(register__n2859) );
  INVx1_ASAP7_75t_R register___U1683 ( .A(register__n2859), .Y(register__n524) );
  OR2x2_ASAP7_75t_R register___U1684 ( .A(register__n370), .B(register__n11580), .Y(register__n1278) );
  NAND4xp25_ASAP7_75t_R register___U1685 ( .A(register__n6713), .B(register__n6711), .C(register__n6825), .D(register__n4720), 
        .Y(register__n370) );
  BUFx6f_ASAP7_75t_R register___U1686 ( .A(register__n12309), .Y(register__n3602) );
  NOR2x1p5_ASAP7_75t_R register___U1687 ( .A(register__n2377), .B(register__n_cell_124812_net160756), .Y(
        n2379) );
  BUFx4_ASAP7_75t_R register___U1688 ( .A(register__net64818), .Y(register__net64788) );
  BUFx4f_ASAP7_75t_R register___U1689 ( .A(register__n12480), .Y(register__n4771) );
  BUFx3_ASAP7_75t_R register___U1690 ( .A(register__n12480), .Y(register__n3704) );
  BUFx12f_ASAP7_75t_R register___U1691 ( .A(register__n3002), .Y(register__n2985) );
  BUFx6f_ASAP7_75t_R register___U1692 ( .A(register__net142400), .Y(register__net64056) );
  INVx2_ASAP7_75t_R register___U1693 ( .A(register__n5480), .Y(register__n9194) );
  INVx6_ASAP7_75t_R register___U1694 ( .A(register__net64790), .Y(register__net64774) );
  INVx1_ASAP7_75t_R register___U1695 ( .A(register__n1303), .Y(register__n1304) );
  OAI22x1_ASAP7_75t_R register___U1696 ( .A1(register__net66310), .A2(register__n7887), .B1(register__n12237), .B2(
        n1687), .Y(read_reg_data_2[17]) );
  BUFx6f_ASAP7_75t_R register___U1697 ( .A(register__n6721), .Y(register__n5181) );
  HB1xp67_ASAP7_75t_R register___U1698 ( .A(register__n4008), .Y(register__n4007) );
  NAND2xp5_ASAP7_75t_R register___U1699 ( .A(register__n1154), .B(register__n1155), .Y(register__n371) );
  BUFx6f_ASAP7_75t_R register___U1700 ( .A(register__net144708), .Y(register__net144463) );
  BUFx6f_ASAP7_75t_R register___U1701 ( .A(register__net144464), .Y(register__net144708) );
  BUFx6f_ASAP7_75t_R register___U1702 ( .A(register__n4270), .Y(register__n3309) );
  INVx2_ASAP7_75t_R register___U1703 ( .A(register__n11826), .Y(register__n11905) );
  OAI22xp33_ASAP7_75t_R register___U1704 ( .A1(register__n12193), .A2(register__n399), .B1(register__n10040), .B2(register__n5641), .Y(register__n372) );
  BUFx4f_ASAP7_75t_R register___U1705 ( .A(register__n7295), .Y(register__n12306) );
  BUFx4f_ASAP7_75t_R register___U1706 ( .A(register__n7296), .Y(register__n3446) );
  INVx2_ASAP7_75t_R register___U1707 ( .A(register__n12306), .Y(register__n12291) );
  AOI22xp33_ASAP7_75t_R register___U1708 ( .A1(register__C6423_net60456), .A2(register__n9503), .B1(
        C6423_net60458), .B2(register__n9445), .Y(register__n11546) );
  AND2x2_ASAP7_75t_R register___U1709 ( .A(register__n7020), .B(register__n7996), .Y(register__C6423_net60458) );
  NOR2xp33_ASAP7_75t_R register___U1710 ( .A(register__C6422_net59832), .B(register__n353), .Y(register__n2494) );
  INVx3_ASAP7_75t_R register___U1711 ( .A(register__n12158), .Y(register__n12147) );
  BUFx6f_ASAP7_75t_R register___U1712 ( .A(register__n3650), .Y(register__n12158) );
  HB1xp67_ASAP7_75t_R register___U1713 ( .A(register__C6423_net61326), .Y(register__net128122) );
  OAI22xp5_ASAP7_75t_R register___U1714 ( .A1(register__n1397), .A2(register__net117656), .B1(register__n1399), .B2(
        n833), .Y(register__n11066) );
  INVxp67_ASAP7_75t_R register___U1715 ( .A(register__C6423_net61348), .Y(register__n631) );
  OAI21xp5_ASAP7_75t_R register___U1716 ( .A1(register__net66310), .A2(register__n2686), .B(register__n2689), .Y(
        read_reg_data_2[15]) );
  BUFx6f_ASAP7_75t_R register___U1717 ( .A(register__n3382), .Y(register__n3380) );
  INVxp33_ASAP7_75t_R register___U1718 ( .A(register__net130175), .Y(register__n373) );
  HB1xp67_ASAP7_75t_R register___U1719 ( .A(register__n13023), .Y(register__n4219) );
  INVx1_ASAP7_75t_R register___U1720 ( .A(register__n12657), .Y(register__n6754) );
  BUFx6f_ASAP7_75t_R register___U1721 ( .A(register__net104685), .Y(register__net137418) );
  BUFx6f_ASAP7_75t_R register___U1722 ( .A(register__n7050), .Y(register__n3938) );
  BUFx3_ASAP7_75t_R register___U1723 ( .A(register__n4033), .Y(register__n3991) );
  CKINVDCx16_ASAP7_75t_R register___U1724 ( .A(register__n11917), .Y(register__n4033) );
  NAND2xp5_ASAP7_75t_R register___U1725 ( .A(register__n8524), .B(register__n59), .Y(register__n412) );
  BUFx2_ASAP7_75t_R register___U1726 ( .A(register__net130175), .Y(register__C6423_net68516) );
  INVx1_ASAP7_75t_R register___U1727 ( .A(register__n13036), .Y(register__n374) );
  BUFx4f_ASAP7_75t_R register___U1728 ( .A(register__n12017), .Y(register__n12004) );
  BUFx12f_ASAP7_75t_R register___U1729 ( .A(register__n11999), .Y(register__n4199) );
  INVx1_ASAP7_75t_R register___U1730 ( .A(register__n12002), .Y(register__n11986) );
  AO22x1_ASAP7_75t_R register___U1731 ( .A1(register__n9718), .A2(register__C6422_net60422), .B1(register__net123857), 
        .B2(register__n10094), .Y(register__n10772) );
  INVxp67_ASAP7_75t_R register___U1732 ( .A(register__n13296), .Y(register__n7276) );
  BUFx2_ASAP7_75t_R register___U1733 ( .A(register__n7706), .Y(register__n8094) );
  INVx4_ASAP7_75t_R register___U1734 ( .A(register__n1139), .Y(register__n1058) );
  INVx2_ASAP7_75t_R register___U1735 ( .A(register__n12493), .Y(register__n1137) );
  INVx1_ASAP7_75t_R register___U1736 ( .A(register__n11520), .Y(register__n376) );
  BUFx6f_ASAP7_75t_R register___U1737 ( .A(register__net66310), .Y(register__net66312) );
  INVx1_ASAP7_75t_R register___U1738 ( .A(register__n10700), .Y(register__n377) );
  NAND2xp67_ASAP7_75t_R register___U1739 ( .A(register__n867), .B(register__n2733), .Y(register__n2687) );
  INVx4_ASAP7_75t_R register___U1740 ( .A(register__n11881), .Y(register__n2016) );
  BUFx6f_ASAP7_75t_R register___U1741 ( .A(register__net131654), .Y(register__n1965) );
  INVx1_ASAP7_75t_R register___U1742 ( .A(register__n13373), .Y(register__n378) );
  NAND2x1p5_ASAP7_75t_R register___U1743 ( .A(register__n149), .B(register__n820), .Y(register__n1872) );
  NAND2x1p5_ASAP7_75t_R register___U1744 ( .A(register__n2402), .B(register__n1284), .Y(register__n754) );
  INVx2_ASAP7_75t_R register___U1745 ( .A(register__C6423_net60460), .Y(register__n711) );
  INVx1_ASAP7_75t_R register___U1746 ( .A(register__n12830), .Y(register__n6726) );
  INVx1_ASAP7_75t_R register___U1747 ( .A(register__n4974), .Y(register__n2928) );
  INVx1_ASAP7_75t_R register___U1748 ( .A(register__n12627), .Y(register__n379) );
  AND3x1_ASAP7_75t_R register___U1749 ( .A(register__n7648), .B(register__n8382), .C(register__n7649), .Y(register__n380) );
  INVx1_ASAP7_75t_R register___U1750 ( .A(register__n6235), .Y(register__n8382) );
  INVx1_ASAP7_75t_R register___U1751 ( .A(register__n12390), .Y(register__n12375) );
  OAI22xp33_ASAP7_75t_R register___U1752 ( .A1(register__n12055), .A2(register__n11876), .B1(register__n9337), .B2(
        n3351), .Y(register__n382) );
  INVx3_ASAP7_75t_R register___U1753 ( .A(register__n9223), .Y(register__n6005) );
  BUFx3_ASAP7_75t_R register___U1754 ( .A(register__net147145), .Y(register__net125384) );
  BUFx6f_ASAP7_75t_R register___U1755 ( .A(register__net125384), .Y(register__net140270) );
  INVx2_ASAP7_75t_R register___U1756 ( .A(register__n6009), .Y(register__n9239) );
  INVx2_ASAP7_75t_R register___U1757 ( .A(register__n10389), .Y(register__n11687) );
  HB1xp67_ASAP7_75t_R register___U1758 ( .A(register__n3450), .Y(register__n3425) );
  BUFx3_ASAP7_75t_R register___U1759 ( .A(register__n12503), .Y(register__n1985) );
  INVx1_ASAP7_75t_R register___U1760 ( .A(register__n12620), .Y(register__n386) );
  AND3x2_ASAP7_75t_R register___U1761 ( .A(register__n572), .B(IF_ID_rs1[2]), .C(register__n11132), .Y(
        n11142) );
  HB1xp67_ASAP7_75t_R register___U1762 ( .A(register__n6498), .Y(register__n6497) );
  INVx2_ASAP7_75t_R register___U1763 ( .A(register__n739), .Y(register__n1036) );
  HB1xp67_ASAP7_75t_R register___U1764 ( .A(register__n3349), .Y(register__n3326) );
  INVx2_ASAP7_75t_R register___U1765 ( .A(register__n277), .Y(register__n2001) );
  INVx1_ASAP7_75t_R register___U1766 ( .A(register__n12940), .Y(register__n390) );
  INVx6_ASAP7_75t_R register___U1767 ( .A(write_data[19]), .Y(register__n12309) );
  INVx1_ASAP7_75t_R register___U1768 ( .A(register__n12960), .Y(register__n391) );
  HB1xp67_ASAP7_75t_R register___U1769 ( .A(register__n12393), .Y(register__n3299) );
  INVxp33_ASAP7_75t_R register___U1770 ( .A(register__n428), .Y(register__n849) );
  NOR2x1p5_ASAP7_75t_R register___U1771 ( .A(register__n2399), .B(register__n2380), .Y(register__n2402) );
  INVx2_ASAP7_75t_R register___U1772 ( .A(register__n4820), .Y(register__n8249) );
  INVx2_ASAP7_75t_R register___U1773 ( .A(register__n12502), .Y(register__n1118) );
  BUFx5_ASAP7_75t_R register___U1774 ( .A(register__n2964), .Y(register__n2963) );
  OAI22xp5_ASAP7_75t_R register___U1775 ( .A1(register__net66302), .A2(register__n7612), .B1(register__n12001), .B2(
        n1687), .Y(read_reg_data_2[2]) );
  BUFx6f_ASAP7_75t_R register___U1776 ( .A(register__net130838), .Y(register__net64060) );
  INVx1_ASAP7_75t_R register___U1777 ( .A(register__n12859), .Y(register__n392) );
  AND2x4_ASAP7_75t_R register___U1778 ( .A(register__net62700), .B(register__n1937), .Y(register__n393) );
  AND2x2_ASAP7_75t_R register___U1779 ( .A(register__n774), .B(register__n2814), .Y(register__n394) );
  NOR2x1p5_ASAP7_75t_R register___U1780 ( .A(register__n393), .B(register__n394), .Y(register__n12859) );
  INVxp33_ASAP7_75t_R register___U1781 ( .A(register__n9515), .Y(register__n774) );
  HB1xp67_ASAP7_75t_R register___U1782 ( .A(register__n2804), .Y(register__n2814) );
  HB1xp67_ASAP7_75t_R register___U1783 ( .A(register__n4662), .Y(register__n4661) );
  INVxp67_ASAP7_75t_R register___U1784 ( .A(register__n3245), .Y(register__n8227) );
  BUFx3_ASAP7_75t_R register___U1785 ( .A(register__n334), .Y(register__net138028) );
  XNOR2x2_ASAP7_75t_R register___U1786 ( .A(register__n154), .B(register__n5441), .Y(register__n12506) );
  AOI22xp33_ASAP7_75t_R register___U1787 ( .A1(register__n12389), .A2(register__n4270), .B1(register__n1052), .B2(register__n1981), .Y(register__n12586) );
  AO22x1_ASAP7_75t_R register___U1788 ( .A1(register__net64788), .A2(register__n5341), .B1(register__n396), .B2(register__n3119), 
        .Y(register__n395) );
  CKINVDCx20_ASAP7_75t_R register___U1789 ( .A(register__net89817), .Y(register__n396) );
  INVx4_ASAP7_75t_R register___U1790 ( .A(register__n3381), .Y(register__n3119) );
  INVx4_ASAP7_75t_R register___U1791 ( .A(register__n3069), .Y(register__n12255) );
  BUFx3_ASAP7_75t_R register___U1792 ( .A(register__n12278), .Y(register__n12277) );
  CKINVDCx20_ASAP7_75t_R register___U1793 ( .A(register__n9437), .Y(register__n397) );
  INVx2_ASAP7_75t_R register___U1794 ( .A(register__n12221), .Y(register__n12204) );
  OAI22xp5_ASAP7_75t_R register___U1795 ( .A1(register__n54), .A2(register__n8645), .B1(register__net61369), .B2(register__n12352), .Y(read_reg_data_1[21]) );
  INVx3_ASAP7_75t_R register___U1796 ( .A(write_data[11]), .Y(register__net64398) );
  INVx2_ASAP7_75t_R register___U1797 ( .A(register__net64352), .Y(register__n456) );
  INVx6_ASAP7_75t_R register___U1798 ( .A(register__net141957), .Y(register__net64352) );
  NOR4xp25_ASAP7_75t_R register___U1799 ( .A(register__n1480), .B(register__n11383), .C(register__n2895), .D(register__n1481), 
        .Y(register__n11365) );
  INVx1_ASAP7_75t_R register___U1800 ( .A(register__n3247), .Y(register__n1481) );
  AND4x1_ASAP7_75t_R register___U1801 ( .A(register__n1437), .B(register__n6748), .C(register__n7263), .D(register__n1319), .Y(
        n11367) );
  AND2x2_ASAP7_75t_R register___U1802 ( .A(register__n10549), .B(register__n10548), .Y(register__n398) );
  AND2x2_ASAP7_75t_R register___U1803 ( .A(register__n1461), .B(register__n398), .Y(register__n7942) );
  INVx5_ASAP7_75t_R register___U1804 ( .A(register__n12486), .Y(register__n399) );
  NOR2xp67_ASAP7_75t_R register___U1805 ( .A(register__n3371), .B(register__n311), .Y(register__n3177) );
  NOR2xp33_ASAP7_75t_R register___U1806 ( .A(register__n12234), .B(register__n338), .Y(register__n400) );
  NOR2x1_ASAP7_75t_R register___U1807 ( .A(register__n9881), .B(register__n343), .Y(register__n401) );
  NOR2xp67_ASAP7_75t_R register___U1808 ( .A(register__n400), .B(register__n401), .Y(register__n12730) );
  BUFx12f_ASAP7_75t_R register___U1809 ( .A(register__net142813), .Y(register__net64886) );
  AND2x2_ASAP7_75t_R register___U1810 ( .A(register__n6199), .B(register__n3130), .Y(register__n402) );
  AND3x1_ASAP7_75t_R register___U1811 ( .A(register__n402), .B(register__n6197), .C(register__n3820), .Y(register__n10590) );
  INVx6_ASAP7_75t_R register___U1812 ( .A(register__n12388), .Y(register__n12376) );
  INVx1_ASAP7_75t_R register___U1813 ( .A(register__n12614), .Y(register__n403) );
  INVxp33_ASAP7_75t_R register___U1814 ( .A(register__n912), .Y(register__n922) );
  HB1xp67_ASAP7_75t_R register___U1815 ( .A(register__n13034), .Y(register__n3580) );
  INVx2_ASAP7_75t_R register___U1816 ( .A(register__net64960), .Y(register__net64928) );
  INVx1_ASAP7_75t_R register___U1817 ( .A(register__n12536), .Y(register__n404) );
  INVx1_ASAP7_75t_R register___U1818 ( .A(register__n11234), .Y(register__n405) );
  INVxp67_ASAP7_75t_R register___U1819 ( .A(register__n2015), .Y(register__net149933) );
  HB1xp67_ASAP7_75t_R register___U1820 ( .A(register__n8095), .Y(register__n7706) );
  INVx3_ASAP7_75t_R register___U1821 ( .A(register__net91939), .Y(register__net64414) );
  OAI22xp33_ASAP7_75t_R register___U1822 ( .A1(register__n1856), .A2(register__n388), .B1(register__n1857), .B2(register__n1336), 
        .Y(register__n10727) );
  OAI22x1_ASAP7_75t_R register___U1823 ( .A1(register__n12373), .A2(register__n2220), .B1(register__n9929), .B2(register__n535), 
        .Y(register__n610) );
  INVx6_ASAP7_75t_R register___U1824 ( .A(register__n3024), .Y(register__n12373) );
  INVx1_ASAP7_75t_R register___U1825 ( .A(register__n13047), .Y(register__n409) );
  INVx1_ASAP7_75t_R register___U1826 ( .A(rs2[1]), .Y(register__n731) );
  NAND2xp33_ASAP7_75t_R register___U1827 ( .A(register__n9849), .B(register__C6422_net60415), .Y(register__n411) );
  NAND2xp33_ASAP7_75t_R register___U1828 ( .A(register__n412), .B(register__n411), .Y(register__n10692) );
  HB1xp67_ASAP7_75t_R register___U1829 ( .A(register__n10299), .Y(register__n8524) );
  BUFx6f_ASAP7_75t_R register___U1830 ( .A(register__n375), .Y(register__C6422_net75149) );
  INVx4_ASAP7_75t_R register___U1831 ( .A(register__C6422_net75149), .Y(register__n_cell_124812_net160756) );
  NOR2xp33_ASAP7_75t_R register___U1832 ( .A(register__n1995), .B(register__n5952), .Y(register__n415) );
  NOR2xp33_ASAP7_75t_R register___U1833 ( .A(register__n1800), .B(register__n6208), .Y(register__n416) );
  NOR3xp33_ASAP7_75t_R register___U1834 ( .A(register__n414), .B(register__n415), .C(register__n416), .Y(register__n11198) );
  HB1xp67_ASAP7_75t_R register___U1835 ( .A(register__n11205), .Y(register__n5952) );
  HB1xp67_ASAP7_75t_R register___U1836 ( .A(register__n11206), .Y(register__n6208) );
  AND2x2_ASAP7_75t_R register___U1837 ( .A(register__n3948), .B(register__n417), .Y(register__n8607) );
  OAI22xp33_ASAP7_75t_R register___U1838 ( .A1(register__n3723), .A2(register__n11859), .B1(register__n10048), .B2(
        n5341), .Y(register__n418) );
  INVx2_ASAP7_75t_R register___U1839 ( .A(register__n7110), .Y(register__n8560) );
  HB1xp67_ASAP7_75t_R register___U1840 ( .A(Reg_data[330]), .Y(register__net103440) );
  INVx2_ASAP7_75t_R register___U1841 ( .A(register__net96598), .Y(register__C6422_net59835) );
  INVx1_ASAP7_75t_R register___U1842 ( .A(register__n12736), .Y(register__n421) );
  INVxp67_ASAP7_75t_R register___U1843 ( .A(register__n475), .Y(register__n4850) );
  INVxp67_ASAP7_75t_R register___U1844 ( .A(register__n12498), .Y(register__n2803) );
  AO22x1_ASAP7_75t_R register___U1845 ( .A1(register__n9744), .A2(register__n3), .B1(register__n10132), .B2(register__n281), .Y(
        n10778) );
  HB1xp67_ASAP7_75t_R register___U1846 ( .A(register__n11386), .Y(register__n7300) );
  AND2x4_ASAP7_75t_R register___U1847 ( .A(register__n11728), .B(register__n441), .Y(register__net122862) );
  INVxp33_ASAP7_75t_R register___U1848 ( .A(register__n1998), .Y(register__net150875) );
  HB1xp67_ASAP7_75t_R register___U1849 ( .A(register__n12619), .Y(register__n4662) );
  OAI22xp33_ASAP7_75t_R register___U1850 ( .A1(register__n12171), .A2(register__n11864), .B1(register__n10140), .B2(
        n5341), .Y(register__n423) );
  OR2x2_ASAP7_75t_R register___U1851 ( .A(register__n652), .B(register__n11726), .Y(register__n651) );
  OR2x6_ASAP7_75t_R register___U1852 ( .A(rs2[3]), .B(rs2[4]), 
        .Y(register__n11726) );
  INVxp33_ASAP7_75t_R register___U1853 ( .A(register__n1439), .Y(register__n1443) );
  INVxp33_ASAP7_75t_R register___U1854 ( .A(register__n1439), .Y(register__n1442) );
  HB1xp67_ASAP7_75t_R register___U1855 ( .A(Reg_data[863]), .Y(register__net103386) );
  HB1xp67_ASAP7_75t_R register___U1856 ( .A(register__C6423_net61304), .Y(register__net111194) );
  HB1xp67_ASAP7_75t_R register___U1857 ( .A(register__net103386), .Y(register__net103385) );
  INVxp67_ASAP7_75t_R register___U1858 ( .A(register__net111194), .Y(register__n543) );
  INVx6_ASAP7_75t_R register___U1859 ( .A(register__net64942), .Y(register__net134981) );
  NAND2xp33_ASAP7_75t_R register___U1860 ( .A(register__n7061), .B(register__n11219), .Y(register__n875) );
  HB1xp67_ASAP7_75t_R register___U1861 ( .A(register__n11220), .Y(register__n7061) );
  AND2x2_ASAP7_75t_R register___U1862 ( .A(register__C6423_net60462), .B(register__n9211), .Y(register__n766) );
  INVxp67_ASAP7_75t_R register___U1863 ( .A(register__n4148), .Y(register__n5371) );
  HB1xp67_ASAP7_75t_R register___U1864 ( .A(register__n4149), .Y(register__n4148) );
  INVxp67_ASAP7_75t_R register___U1865 ( .A(register__n1013), .Y(register__n1014) );
  NOR3x1_ASAP7_75t_R register___U1866 ( .A(register__n5810), .B(register__n8746), .C(register__n8744), .Y(register__n424) );
  NOR2xp67_ASAP7_75t_R register___U1867 ( .A(register__n817), .B(register__C6423_net60882), .Y(register__n497) );
  HB1xp67_ASAP7_75t_R register___U1868 ( .A(register__n7652), .Y(register__n3111) );
  BUFx12f_ASAP7_75t_R register___U1869 ( .A(register__net141991), .Y(register__net141459) );
  NAND2xp67_ASAP7_75t_R register___U1870 ( .A(register__n756), .B(register__n11174), .Y(register__n425) );
  NOR3x1_ASAP7_75t_R register___U1871 ( .A(register__n5414), .B(register__n5409), .C(register__n5248), .Y(register__n756) );
  BUFx3_ASAP7_75t_R register___U1872 ( .A(register__n3512), .Y(register__n8247) );
  HB1xp67_ASAP7_75t_R register___U1873 ( .A(register__n13334), .Y(register__n5014) );
  HB1xp67_ASAP7_75t_R register___U1874 ( .A(register__n13305), .Y(register__n4874) );
  NOR2xp33_ASAP7_75t_R register___U1875 ( .A(register__n1995), .B(register__n9157), .Y(register__n2753) );
  INVx1_ASAP7_75t_R register___U1876 ( .A(register__n12542), .Y(register__n426) );
  INVx2_ASAP7_75t_R register___U1877 ( .A(register__n456), .Y(register__net64344) );
  AND3x2_ASAP7_75t_R register___U1878 ( .A(register__n7067), .B(register__n29), .C(register__n7068), .Y(register__n427) );
  AND2x2_ASAP7_75t_R register___U1879 ( .A(register__n7069), .B(register__n427), .Y(register__n10613) );
  HB1xp67_ASAP7_75t_R register___U1880 ( .A(register__n3183), .Y(register__n3182) );
  HB1xp67_ASAP7_75t_R register___U1881 ( .A(register__n11725), .Y(register__n3183) );
  CKINVDCx10_ASAP7_75t_R register___U1882 ( .A(register__net128430), .Y(register__net64942) );
  INVxp33_ASAP7_75t_R register___U1883 ( .A(register__n2015), .Y(register__net149938) );
  INVxp33_ASAP7_75t_R register___U1884 ( .A(register__n2015), .Y(register__net149939) );
  HB1xp67_ASAP7_75t_R register___U1885 ( .A(IF_ID_rs1[1]), .Y(register__n428) );
  HB1xp67_ASAP7_75t_R register___U1886 ( .A(IF_ID_rs1[1]), .Y(register__n429) );
  HB1xp67_ASAP7_75t_R register___U1887 ( .A(IF_ID_rs1[1]), .Y(register__n1476) );
  NAND2xp5_ASAP7_75t_R register___U1888 ( .A(register__n8202), .B(register__n834), .Y(register__n863) );
  INVxp67_ASAP7_75t_R register___U1889 ( .A(register__n3554), .Y(register__n4184) );
  HB1xp67_ASAP7_75t_R register___U1890 ( .A(register__n3555), .Y(register__n3554) );
  HB1xp67_ASAP7_75t_R register___U1891 ( .A(register__n12812), .Y(register__n3555) );
  HB1xp67_ASAP7_75t_R register___U1892 ( .A(register__n3598), .Y(register__n3453) );
  INVxp67_ASAP7_75t_R register___U1893 ( .A(register__n5803), .Y(register__n8300) );
  BUFx3_ASAP7_75t_R register___U1894 ( .A(register__n11874), .Y(register__n11755) );
  OR2x6_ASAP7_75t_R register___U1895 ( .A(register__n2167), .B(register__n12491), .Y(register__n7633) );
  HB1xp67_ASAP7_75t_R register___U1896 ( .A(register__n6801), .Y(register__n3444) );
  HB1xp67_ASAP7_75t_R register___U1897 ( .A(WB_rd[3]), .Y(register__n4264) );
  INVx1_ASAP7_75t_R register___U1898 ( .A(register__n729), .Y(register__n1489) );
  HB1xp67_ASAP7_75t_R register___U1899 ( .A(register__n5426), .Y(register__n5425) );
  BUFx3_ASAP7_75t_R register___U1900 ( .A(register__n3473), .Y(register__n6301) );
  INVx1_ASAP7_75t_R register___U1901 ( .A(register__n12687), .Y(register__n431) );
  NAND2xp33_ASAP7_75t_R register___U1902 ( .A(register__n1110), .B(register__n195), .Y(register__n433) );
  AND2x2_ASAP7_75t_R register___U1903 ( .A(register__n432), .B(register__n433), .Y(register__n12687) );
  BUFx6f_ASAP7_75t_R register___U1904 ( .A(register__n3389), .Y(register__n11899) );
  INVxp33_ASAP7_75t_R register___U1905 ( .A(register__n8757), .Y(register__n1110) );
  BUFx12f_ASAP7_75t_R register___U1906 ( .A(register__n5503), .Y(register__n5501) );
  INVxp33_ASAP7_75t_R register___U1907 ( .A(register__net94400), .Y(register__n435) );
  HB1xp67_ASAP7_75t_R register___U1908 ( .A(register__net94400), .Y(register__n436) );
  BUFx6f_ASAP7_75t_R register___U1909 ( .A(register__n515), .Y(register__C6423_net68914) );
  BUFx6f_ASAP7_75t_R register___U1910 ( .A(register__C6423_net68914), .Y(register__net94399) );
  INVx1_ASAP7_75t_R register___U1911 ( .A(register__n13039), .Y(register__n438) );
  AO22x1_ASAP7_75t_R register___U1912 ( .A1(register__n10434), .A2(register__net91683), .B1(register__n10421), .B2(
        n1347), .Y(register__n10688) );
  BUFx12f_ASAP7_75t_R register___U1913 ( .A(register__net142807), .Y(register__net62700) );
  BUFx12f_ASAP7_75t_R register___U1914 ( .A(register__n12473), .Y(register__n3348) );
  INVx1_ASAP7_75t_R register___U1915 ( .A(register__n12997), .Y(register__n439) );
  INVxp67_ASAP7_75t_R register___U1916 ( .A(register__n12919), .Y(register__n6135) );
  INVx1_ASAP7_75t_R register___U1917 ( .A(register__n429), .Y(register__n729) );
  OAI22xp33_ASAP7_75t_R register___U1918 ( .A1(register__n12457), .A2(register__n957), .B1(register__n9315), .B2(register__n958), 
        .Y(register__n440) );
  BUFx2_ASAP7_75t_R register___U1919 ( .A(register__n8370), .Y(register__n8978) );
  AND2x2_ASAP7_75t_R register___U1920 ( .A(register__n9389), .B(register__n1128), .Y(register__n5951) );
  NAND2xp5_ASAP7_75t_R register___U1921 ( .A(register__n12503), .B(register__n5951), .Y(register__n475) );
  INVx1_ASAP7_75t_R register___U1922 ( .A(register__n11475), .Y(register__n8284) );
  HB1xp67_ASAP7_75t_R register___U1923 ( .A(register__n12729), .Y(register__n3286) );
  OAI22xp5_ASAP7_75t_R register___U1924 ( .A1(register__net66320), .A2(register__n4179), .B1(register__n12466), .B2(
        n1687), .Y(read_reg_data_2[30]) );
  INVxp67_ASAP7_75t_R register___U1925 ( .A(register__n1606), .Y(register__n12845) );
  AND3x2_ASAP7_75t_R register___U1926 ( .A(register__n3642), .B(register__n3943), .C(register__n3641), .Y(register__n442) );
  AND2x2_ASAP7_75t_R register___U1927 ( .A(register__n3042), .B(register__n442), .Y(register__n10757) );
  INVx1_ASAP7_75t_R register___U1928 ( .A(register__n3039), .Y(register__n3641) );
  INVx2_ASAP7_75t_R register___U1929 ( .A(register__net88572), .Y(register__net117656) );
  INVxp67_ASAP7_75t_R register___U1930 ( .A(register__n1773), .Y(register__n1381) );
  INVxp33_ASAP7_75t_R register___U1931 ( .A(register__n109), .Y(register__n567) );
  INVxp33_ASAP7_75t_R register___U1932 ( .A(register__n109), .Y(register__n1379) );
  AND2x4_ASAP7_75t_R register___U1933 ( .A(register__n565), .B(register__n8752), .Y(register__n443) );
  BUFx3_ASAP7_75t_R register___U1934 ( .A(register__n10801), .Y(register__n8638) );
  NOR2xp67_ASAP7_75t_R register___U1935 ( .A(register__n9199), .B(register__n27), .Y(register__n1021) );
  AND2x4_ASAP7_75t_R register___U1936 ( .A(IF_ID_rs1[2]), .B(register__n11136), .Y(register__n11135) );
  INVx1_ASAP7_75t_R register___U1937 ( .A(register__n13299), .Y(register__n444) );
  INVx4_ASAP7_75t_R register___U1938 ( .A(register__n12249), .Y(register__n781) );
  INVxp33_ASAP7_75t_R register___U1939 ( .A(register__n733), .Y(register__n12227) );
  NOR2xp33_ASAP7_75t_R register___U1940 ( .A(register__net64942), .B(register__n105), .Y(register__n2314) );
  INVx3_ASAP7_75t_R register___U1941 ( .A(register__n12239), .Y(register__n12226) );
  OAI22xp33_ASAP7_75t_R register___U1942 ( .A1(register__n11926), .A2(register__n889), .B1(register__n9411), .B2(register__n905), 
        .Y(register__n445) );
  HB1xp67_ASAP7_75t_R register___U1943 ( .A(register__n11421), .Y(register__n5426) );
  AO22x1_ASAP7_75t_R register___U1944 ( .A1(register__n8805), .A2(register__net117658), .B1(register__n7337), .B2(register__n839), 
        .Y(register__n10871) );
  AO22x1_ASAP7_75t_R register___U1945 ( .A1(register__n9272), .A2(register__C6422_net60408), .B1(register__n10237), 
        .B2(register__n837), .Y(register__n10894) );
  AO22x1_ASAP7_75t_R register___U1946 ( .A1(register__net93468), .A2(register__C6422_net60408), .B1(register__net93408), 
        .B2(register__n841), .Y(register__n11085) );
  INVxp67_ASAP7_75t_R register___U1947 ( .A(register__n4527), .Y(register__n6185) );
  INVxp67_ASAP7_75t_R register___U1948 ( .A(register__n5091), .Y(register__n7043) );
  AO22x1_ASAP7_75t_R register___U1949 ( .A1(register__n4290), .A2(register__n1697), .B1(register__n446), .B2(register__n1714), 
        .Y(register__n1401) );
  CKINVDCx20_ASAP7_75t_R register___U1950 ( .A(register__n8803), .Y(register__n446) );
  OAI22xp33_ASAP7_75t_R register___U1951 ( .A1(register__n11926), .A2(register__n951), .B1(register__n9658), .B2(register__n958), 
        .Y(register__n447) );
  NOR2xp33_ASAP7_75t_R register___U1952 ( .A(register__n2217), .B(register__n2216), .Y(register__n3994) );
  OAI22xp33_ASAP7_75t_R register___U1953 ( .A1(register__n53), .A2(register__n3994), .B1(register__net61369), .B2(
        net64360), .Y(read_reg_data_1[11]) );
  INVx1_ASAP7_75t_R register___U1954 ( .A(register__n1299), .Y(register__n448) );
  INVxp33_ASAP7_75t_R register___U1955 ( .A(register__n1299), .Y(register__n6466) );
  OAI22xp5_ASAP7_75t_R register___U1956 ( .A1(register__n53), .A2(register__n8586), .B1(register__net61369), .B2(
        net64974), .Y(read_reg_data_1[4]) );
  NAND2xp33_ASAP7_75t_R register___U1957 ( .A(register__n9347), .B(register__net117657), .Y(register__n1514) );
  INVxp67_ASAP7_75t_R register___U1958 ( .A(register__n11944), .Y(register__n11930) );
  INVxp67_ASAP7_75t_R register___U1959 ( .A(register__n11942), .Y(register__n11929) );
  AO22x1_ASAP7_75t_R register___U1960 ( .A1(register__net138525), .A2(register__n2020), .B1(register__n450), .B2(register__n451), 
        .Y(register__n449) );
  CKINVDCx20_ASAP7_75t_R register___U1961 ( .A(register__net89717), .Y(register__n450) );
  INVx13_ASAP7_75t_R register___U1962 ( .A(register__n11850), .Y(register__n451) );
  INVxp33_ASAP7_75t_R register___U1963 ( .A(register__n4816), .Y(register__n11931) );
  BUFx4f_ASAP7_75t_R register___U1964 ( .A(register__net141508), .Y(register__net122410) );
  BUFx4f_ASAP7_75t_R register___U1965 ( .A(register__net122410), .Y(register__net140640) );
  HB1xp67_ASAP7_75t_R register___U1966 ( .A(register__n7656), .Y(register__n3306) );
  HB1xp67_ASAP7_75t_R register___U1967 ( .A(register__n12500), .Y(register__n7656) );
  AOI21xp5_ASAP7_75t_R register___U1968 ( .A1(register__n2000), .A2(register__net89585), .B(register__n452), .Y(register__n546)
         );
  AO21x1_ASAP7_75t_R register___U1969 ( .A1(register__C6423_net68914), .A2(register__net89601), .B(register__n2601), 
        .Y(register__n452) );
  INVx2_ASAP7_75t_R register___U1970 ( .A(register__n277), .Y(register__n2000) );
  BUFx3_ASAP7_75t_R register___U1971 ( .A(register__net105786), .Y(register__net89585) );
  INVx2_ASAP7_75t_R register___U1972 ( .A(register__n11939), .Y(register__n11935) );
  INVxp67_ASAP7_75t_R register___U1973 ( .A(register__n5759), .Y(register__n8655) );
  INVxp67_ASAP7_75t_R register___U1974 ( .A(register__C6423_net74857), .Y(register__n453) );
  HB1xp67_ASAP7_75t_R register___U1975 ( .A(register__net147378), .Y(register__net145304) );
  NOR3x1_ASAP7_75t_R register___U1976 ( .A(register__n6005), .B(register__n9224), .C(register__n9222), .Y(register__n455) );
  BUFx12f_ASAP7_75t_R register___U1977 ( .A(register__n2844), .Y(register__n11780) );
  NAND3xp33_ASAP7_75t_R register___U1978 ( .A(register__n10568), .B(register__n6453), .C(register__n10569), .Y(register__n1013)
         );
  NAND2x1p5_ASAP7_75t_R register___U1979 ( .A(register__n546), .B(register__n547), .Y(register__n537) );
  HB1xp67_ASAP7_75t_R register___U1980 ( .A(register__n8979), .Y(register__n8370) );
  BUFx12f_ASAP7_75t_R register___U1981 ( .A(register__n11888), .Y(register__n5838) );
  AO22x1_ASAP7_75t_R register___U1982 ( .A1(register__n9895), .A2(register__n38), .B1(register__n10153), .B2(
        C6422_net60443), .Y(register__n11074) );
  AO22x1_ASAP7_75t_R register___U1983 ( .A1(register__n9634), .A2(register__C6422_net60445), .B1(register__n7478), .B2(
        C6422_net60443), .Y(register__n10543) );
  AO22x1_ASAP7_75t_R register___U1984 ( .A1(register__n9282), .A2(register__n77), .B1(register__n10152), .B2(register__net108158), 
        .Y(register__n10776) );
  INVx2_ASAP7_75t_R register___U1985 ( .A(register__n2998), .Y(register__n6448) );
  INVx1_ASAP7_75t_R register___U1986 ( .A(write_data[30]), .Y(register__n12482) );
  BUFx6f_ASAP7_75t_R register___U1987 ( .A(register__n11782), .Y(register__n457) );
  BUFx4f_ASAP7_75t_R register___U1988 ( .A(register__n11782), .Y(register__n458) );
  INVx2_ASAP7_75t_R register___U1989 ( .A(register__n12496), .Y(register__n460) );
  INVx2_ASAP7_75t_R register___U1990 ( .A(register__n457), .Y(register__n463) );
  INVx2_ASAP7_75t_R register___U1991 ( .A(register__n457), .Y(register__n464) );
  INVx2_ASAP7_75t_R register___U1992 ( .A(register__n457), .Y(register__n465) );
  INVx2_ASAP7_75t_R register___U1993 ( .A(register__n457), .Y(register__n466) );
  INVx2_ASAP7_75t_R register___U1994 ( .A(register__n457), .Y(register__n467) );
  INVx2_ASAP7_75t_R register___U1995 ( .A(register__n457), .Y(register__n468) );
  INVx2_ASAP7_75t_R register___U1996 ( .A(register__n458), .Y(register__n469) );
  INVx2_ASAP7_75t_R register___U1997 ( .A(register__n458), .Y(register__n470) );
  INVx1_ASAP7_75t_R register___U1998 ( .A(register__n458), .Y(register__n471) );
  INVx1_ASAP7_75t_R register___U1999 ( .A(register__n458), .Y(register__n472) );
  INVx1_ASAP7_75t_R register___U2000 ( .A(register__n458), .Y(register__n473) );
  INVx1_ASAP7_75t_R register___U2001 ( .A(register__n458), .Y(register__n474) );
  INVx4_ASAP7_75t_R register___U2002 ( .A(register__n3652), .Y(register__n11782) );
  BUFx2_ASAP7_75t_R register___U2003 ( .A(register__n12496), .Y(register__n3652) );
  INVxp67_ASAP7_75t_R register___U2004 ( .A(register__n12591), .Y(register__n6729) );
  BUFx6f_ASAP7_75t_R register___U2005 ( .A(register__n3344), .Y(register__n11781) );
  BUFx2_ASAP7_75t_R register___U2006 ( .A(register__n3438), .Y(register__n3437) );
  BUFx6f_ASAP7_75t_R register___U2007 ( .A(register__n11869), .Y(register__n3438) );
  AO22x1_ASAP7_75t_R register___U2008 ( .A1(register__n12333), .A2(register__n1603), .B1(register__n477), .B2(register__n11816), 
        .Y(register__n476) );
  CKINVDCx20_ASAP7_75t_R register___U2009 ( .A(register__n9447), .Y(register__n477) );
  NAND2x1p5_ASAP7_75t_R register___U2010 ( .A(register__net62704), .B(register__n5548), .Y(register__n1087) );
  INVxp33_ASAP7_75t_R register___U2011 ( .A(register__n1951), .Y(register__n976) );
  INVx3_ASAP7_75t_R register___U2012 ( .A(register__n2813), .Y(register__n1937) );
  OAI21xp33_ASAP7_75t_R register___U2013 ( .A1(register__net107791), .A2(register__n66), .B(register__n2348), .Y(register__n2347)
         );
  HB1xp67_ASAP7_75t_R register___U2014 ( .A(register__n12845), .Y(register__n5091) );
  AO22x1_ASAP7_75t_R register___U2015 ( .A1(register__net140427), .A2(register__C6423_net61340), .B1(
        net110205), .B2(register__C6423_net69198), .Y(register__n11271) );
  BUFx3_ASAP7_75t_R register___U2016 ( .A(register__n3546), .Y(register__n3673) );
  HB1xp67_ASAP7_75t_R register___U2017 ( .A(register__n13295), .Y(register__n4872) );
  INVxp67_ASAP7_75t_R register___U2018 ( .A(register__n531), .Y(register__n13295) );
  AO22x1_ASAP7_75t_R register___U2019 ( .A1(register__n3265), .A2(register__n5341), .B1(register__n532), .B2(register__n399), .Y(
        n531) );
  INVxp67_ASAP7_75t_R register___U2020 ( .A(register__n596), .Y(register__n1039) );
  HB1xp67_ASAP7_75t_R register___U2021 ( .A(register__n12513), .Y(register__n6761) );
  INVx1_ASAP7_75t_R register___U2022 ( .A(register__n1039), .Y(register__n716) );
  BUFx6f_ASAP7_75t_R register___U2023 ( .A(register__n667), .Y(register__net127751) );
  NOR3x1_ASAP7_75t_R register___U2024 ( .A(register__n5124), .B(register__n7673), .C(register__n7672), .Y(register__n479) );
  AND2x2_ASAP7_75t_R register___U2025 ( .A(register__C6423_net60460), .B(register__n9463), .Y(register__n765) );
  AND2x4_ASAP7_75t_R register___U2026 ( .A(register__n11728), .B(register__n740), .Y(register__C6423_net60460) );
  CKINVDCx20_ASAP7_75t_R register___U2027 ( .A(register__n9889), .Y(register__n480) );
  CKINVDCx5p33_ASAP7_75t_R register___U2028 ( .A(register__n12242), .Y(register__n12230) );
  INVx5_ASAP7_75t_R register___U2029 ( .A(register__n1411), .Y(register__n1417) );
  BUFx4f_ASAP7_75t_R register___U2030 ( .A(register__net141449), .Y(register__net144154) );
  HB1xp67_ASAP7_75t_R register___U2031 ( .A(register__n7592), .Y(register__n12411) );
  INVx6_ASAP7_75t_R register___U2032 ( .A(register__n12405), .Y(register__n7592) );
  AND3x1_ASAP7_75t_R register___U2033 ( .A(register__n483), .B(register__n11175), .C(register__n424), .Y(register__n8338) );
  BUFx2_ASAP7_75t_R register___U2034 ( .A(register__n11948), .Y(register__n11944) );
  BUFx6f_ASAP7_75t_R register___U2035 ( .A(register__n3535), .Y(register__n3534) );
  INVx1_ASAP7_75t_R register___U2036 ( .A(register__n12962), .Y(register__n484) );
  INVxp67_ASAP7_75t_R register___U2037 ( .A(register__n1098), .Y(register__n485) );
  INVx3_ASAP7_75t_R register___U2038 ( .A(register__n3478), .Y(register__n1098) );
  HB1xp67_ASAP7_75t_R register___U2039 ( .A(register__n12738), .Y(register__n3616) );
  BUFx2_ASAP7_75t_R register___U2040 ( .A(register__n4283), .Y(register__n12103) );
  BUFx2_ASAP7_75t_R register___U2041 ( .A(register__n4283), .Y(register__n12104) );
  AO22x1_ASAP7_75t_R register___U2042 ( .A1(register__n8538), .A2(register__n883), .B1(register__n7561), .B2(register__net122862), 
        .Y(register__n11463) );
  NOR2xp67_ASAP7_75t_R register___U2043 ( .A(register__n5051), .B(register__n32), .Y(register__n11080) );
  HB1xp67_ASAP7_75t_R register___U2044 ( .A(register__n11088), .Y(register__n3147) );
  NOR2x1_ASAP7_75t_R register___U2045 ( .A(register__n2705), .B(register__n_cell_125217_net175364), .Y(register__n2706)
         );
  INVxp67_ASAP7_75t_R register___U2046 ( .A(register__n10910), .Y(register__n486) );
  BUFx2_ASAP7_75t_R register___U2047 ( .A(register__n12191), .Y(register__n12190) );
  INVx2_ASAP7_75t_R register___U2048 ( .A(write_data[14]), .Y(register__n12191) );
  HB1xp67_ASAP7_75t_R register___U2049 ( .A(Reg_data[71]), .Y(register__n8979) );
  BUFx6f_ASAP7_75t_R register___U2050 ( .A(register__n9514), .Y(register__n8981) );
  INVx1_ASAP7_75t_R register___U2051 ( .A(register__n12905), .Y(register__n487) );
  AO22x1_ASAP7_75t_R register___U2052 ( .A1(register__n9625), .A2(register__n38), .B1(register__n10088), .B2(register__n369), .Y(
        n10879) );
  NOR2xp33_ASAP7_75t_R register___U2053 ( .A(register__C6423_net61245), .B(register__n1987), .Y(register__n2533) );
  HB1xp67_ASAP7_75t_R register___U2054 ( .A(register__n11176), .Y(register__n5809) );
  HB1xp67_ASAP7_75t_R register___U2055 ( .A(register__n12788), .Y(register__n4532) );
  INVx4_ASAP7_75t_R register___U2056 ( .A(register__n12180), .Y(register__n12168) );
  OR2x6_ASAP7_75t_R register___U2057 ( .A(register__n1036), .B(register__n2739), .Y(register__n488) );
  AO22x1_ASAP7_75t_R register___U2058 ( .A1(register__net138525), .A2(register__n490), .B1(register__n491), .B2(register__n492), 
        .Y(register__n489) );
  CKINVDCx20_ASAP7_75t_R register___U2059 ( .A(register__n11730), .Y(register__n490) );
  CKINVDCx20_ASAP7_75t_R register___U2060 ( .A(register__net88893), .Y(register__n491) );
  CKINVDCx20_ASAP7_75t_R register___U2061 ( .A(register__n1164), .Y(register__n492) );
  INVx4_ASAP7_75t_R register___U2062 ( .A(write_data[2]), .Y(register__n12017) );
  INVx2_ASAP7_75t_R register___U2063 ( .A(register__n4122), .Y(register__n1594) );
  INVx1_ASAP7_75t_R register___U2064 ( .A(register__n11263), .Y(register__n493) );
  INVx6_ASAP7_75t_R register___U2065 ( .A(register__net64062), .Y(register__net142401) );
  INVxp67_ASAP7_75t_R register___U2066 ( .A(register__n4395), .Y(register__n6753) );
  INVxp67_ASAP7_75t_R register___U2067 ( .A(register__n12405), .Y(register__n1249) );
  BUFx4f_ASAP7_75t_R register___U2068 ( .A(register__C6423_net69526), .Y(register__net110413) );
  BUFx6f_ASAP7_75t_R register___U2069 ( .A(register__n3350), .Y(register__n5531) );
  INVxp33_ASAP7_75t_R register___U2070 ( .A(register__n1101), .Y(register__n13084) );
  HB1xp67_ASAP7_75t_R register___U2071 ( .A(register__n13072), .Y(register__n6498) );
  AO22x1_ASAP7_75t_R register___U2072 ( .A1(register__n11942), .A2(register__n4268), .B1(register__n495), .B2(register__n594), 
        .Y(register__n494) );
  CKINVDCx20_ASAP7_75t_R register___U2073 ( .A(register__n9700), .Y(register__n495) );
  NAND2xp5_ASAP7_75t_R register___U2074 ( .A(register__n328), .B(register__n820), .Y(register__n1133) );
  BUFx3_ASAP7_75t_R register___U2075 ( .A(register__n2840), .Y(register__n3560) );
  NOR2xp33_ASAP7_75t_R register___U2076 ( .A(register__n2002), .B(register__net118829), .Y(register__n496) );
  NOR2xp33_ASAP7_75t_R register___U2077 ( .A(register__net106712), .B(register__net112580), .Y(register__n498) );
  NOR3xp33_ASAP7_75t_R register___U2078 ( .A(register__n496), .B(register__n497), .C(register__n498), .Y(register__n10803) );
  INVx2_ASAP7_75t_R register___U2079 ( .A(register__net91307), .Y(register__C6423_net60882) );
  HB1xp67_ASAP7_75t_R register___U2080 ( .A(register__C6422_net59965), .Y(register__net106712) );
  BUFx6f_ASAP7_75t_R register___U2081 ( .A(register__n3600), .Y(register__n8246) );
  HB1xp67_ASAP7_75t_R register___U2082 ( .A(register__net129787), .Y(register__C6423_net69274) );
  AND2x4_ASAP7_75t_R register___U2083 ( .A(register__n877), .B(register__n739), .Y(register__net122313) );
  NAND2xp5_ASAP7_75t_R register___U2085 ( .A(register__n2185), .B(register__n2186), .Y(register__n2188) );
  BUFx6f_ASAP7_75t_R register___U2086 ( .A(register__n5349), .Y(register__n3516) );
  HB1xp67_ASAP7_75t_R register___U2087 ( .A(register__n5804), .Y(register__n5803) );
  HB1xp67_ASAP7_75t_R register___U2088 ( .A(register__n12108), .Y(register__n12107) );
  INVx6_ASAP7_75t_R register___U2089 ( .A(register__n11776), .Y(register__n11877) );
  BUFx3_ASAP7_75t_R register___U2090 ( .A(register__n11748), .Y(register__n11745) );
  OAI22xp33_ASAP7_75t_R register___U2091 ( .A1(register__n11923), .A2(register__n1698), .B1(register__n10016), .B2(
        n1694), .Y(register__n499) );
  OAI22xp5_ASAP7_75t_R register___U2092 ( .A1(register__n53), .A2(register__n8273), .B1(register__net61369), .B2(register__n12065), .Y(read_reg_data_1[8]) );
  NOR2x2_ASAP7_75t_R register___U2093 ( .A(register__C6422_net59731), .B(register__net130087), .Y(register__n2373) );
  INVx2_ASAP7_75t_R register___U2094 ( .A(register__n7020), .Y(register__n1335) );
  INVx2_ASAP7_75t_R register___U2095 ( .A(register__C6423_net60460), .Y(register__n713) );
  HB1xp67_ASAP7_75t_R register___U2096 ( .A(register__n12532), .Y(register__n5750) );
  BUFx12f_ASAP7_75t_R register___U2097 ( .A(register__n4198), .Y(register__n3383) );
  HB1xp67_ASAP7_75t_R register___U2098 ( .A(register__net147584), .Y(register__net147822) );
  BUFx2_ASAP7_75t_R register___U2099 ( .A(register__net147822), .Y(register__net147907) );
  AO22x1_ASAP7_75t_R register___U2100 ( .A1(register__n9278), .A2(register__n77), .B1(register__n9931), .B2(register__n75), .Y(
        n10926) );
  AO22x1_ASAP7_75t_R register___U2101 ( .A1(register__net93713), .A2(register__n77), .B1(register__net89641), .B2(register__n75), 
        .Y(register__n10815) );
  AO22x1_ASAP7_75t_R register___U2102 ( .A1(register__n9913), .A2(register__n77), .B1(register__n10216), .B2(register__n75), .Y(
        n11118) );
  AO22x1_ASAP7_75t_R register___U2103 ( .A1(register__n6980), .A2(register__n77), .B1(register__n10218), .B2(
        C6422_net60437), .Y(register__n10799) );
  AO22x1_ASAP7_75t_R register___U2104 ( .A1(register__n6893), .A2(register__n77), .B1(register__n9323), .B2(
        C6422_net60437), .Y(register__n10836) );
  AO22x1_ASAP7_75t_R register___U2105 ( .A1(register__n9292), .A2(register__n768), .B1(register__n9939), .B2(
        C6422_net60437), .Y(register__n10585) );
  AOI22xp33_ASAP7_75t_R register___U2106 ( .A1(register__net64698), .A2(register__n2816), .B1(register__n9148), .B2(
        n2810), .Y(register__n12880) );
  BUFx6f_ASAP7_75t_R register___U2107 ( .A(register__n12419), .Y(register__n12416) );
  INVx1_ASAP7_75t_R register___U2108 ( .A(register__n12419), .Y(register__n12404) );
  HB1xp67_ASAP7_75t_R register___U2109 ( .A(register__n373), .Y(register__net114704) );
  INVx1_ASAP7_75t_R register___U2110 ( .A(register__n13147), .Y(register__n502) );
  NAND2xp33_ASAP7_75t_R register___U2111 ( .A(register__n11937), .B(register__n3334), .Y(register__n503) );
  NAND2xp33_ASAP7_75t_R register___U2112 ( .A(register__n1265), .B(register__n1755), .Y(register__n504) );
  AND2x2_ASAP7_75t_R register___U2113 ( .A(register__n503), .B(register__n504), .Y(register__n13147) );
  BUFx6f_ASAP7_75t_R register___U2114 ( .A(register__n3594), .Y(register__n11937) );
  INVxp33_ASAP7_75t_R register___U2115 ( .A(register__n9696), .Y(register__n1265) );
  NOR2xp67_ASAP7_75t_R register___U2116 ( .A(register__n857), .B(register__n858), .Y(register__n505) );
  NOR2x1_ASAP7_75t_R register___U2117 ( .A(register__n856), .B(register__n506), .Y(register__n7668) );
  INVx1_ASAP7_75t_R register___U2118 ( .A(register__n505), .Y(register__n506) );
  NOR2xp33_ASAP7_75t_R register___U2119 ( .A(register__net127626), .B(register__C6422_net59703), .Y(register__n856) );
  INVx1_ASAP7_75t_R register___U2120 ( .A(register__n1160), .Y(register__net100543) );
  BUFx6f_ASAP7_75t_R register___U2121 ( .A(register__n775), .Y(register__net64458) );
  INVxp33_ASAP7_75t_R register___U2122 ( .A(register__net147583), .Y(register__n1160) );
  AND2x4_ASAP7_75t_R register___U2123 ( .A(register__n11719), .B(register__n11728), .Y(register__C6423_net61331) );
  INVxp67_ASAP7_75t_R register___U2124 ( .A(register__n8301), .Y(register__n5805) );
  HB1xp67_ASAP7_75t_R register___U2125 ( .A(register__n11521), .Y(register__n8301) );
  INVx4_ASAP7_75t_R register___U2126 ( .A(register__net64446), .Y(register__net64422) );
  INVx1_ASAP7_75t_R register___U2127 ( .A(register__n12589), .Y(register__n508) );
  INVx1_ASAP7_75t_R register___U2128 ( .A(WB_rd[4]), .Y(register__n5247) );
  INVxp67_ASAP7_75t_R register___U2129 ( .A(register__n4105), .Y(register__n6751) );
  AO22x1_ASAP7_75t_R register___U2130 ( .A1(register__n9650), .A2(register__n1909), .B1(register__n9977), .B2(register__n381), 
        .Y(register__n10632) );
  INVx2_ASAP7_75t_R register___U2131 ( .A(WB_rd[2]), .Y(register__n12489) );
  INVx1_ASAP7_75t_R register___U2132 ( .A(register__n12966), .Y(register__n510) );
  AND4x1_ASAP7_75t_R register___U2133 ( .A(register__n7063), .B(register__n7062), .C(register__n8255), .D(register__n1340), .Y(
        n11220) );
  INVx1_ASAP7_75t_R register___U2134 ( .A(register__C6423_net61317), .Y(register__n1441) );
  INVx3_ASAP7_75t_R register___U2135 ( .A(register__n3343), .Y(register__n3344) );
  INVx4_ASAP7_75t_R register___U2136 ( .A(register__n10517), .Y(register__n3343) );
  INVx3_ASAP7_75t_R register___U2137 ( .A(register__n3449), .Y(register__n12457) );
  OAI22xp33_ASAP7_75t_R register___U2138 ( .A1(register__n11923), .A2(register__n11868), .B1(register__n10030), .B2(
        n3560), .Y(register__n511) );
  NOR2xp67_ASAP7_75t_R register___U2139 ( .A(register__n1994), .B(register__net109872), .Y(register__n1033) );
  BUFx6f_ASAP7_75t_R register___U2140 ( .A(register__net100798), .Y(register__net62698) );
  BUFx6f_ASAP7_75t_R register___U2141 ( .A(register__net100799), .Y(register__net100798) );
  AO22x1_ASAP7_75t_R register___U2142 ( .A1(register__n12183), .A2(register__n4851), .B1(register__n513), .B2(register__n1848), 
        .Y(register__n512) );
  CKINVDCx20_ASAP7_75t_R register___U2143 ( .A(register__n9557), .Y(register__n513) );
  INVx1_ASAP7_75t_R register___U2144 ( .A(register__n4851), .Y(register__n698) );
  HB1xp67_ASAP7_75t_R register___U2145 ( .A(register__n12798), .Y(register__n4504) );
  INVx3_ASAP7_75t_R register___U2146 ( .A(register__n1524), .Y(register__n1984) );
  AND2x4_ASAP7_75t_R register___U2147 ( .A(register__n3407), .B(register__n1985), .Y(register__n4270) );
  HB1xp67_ASAP7_75t_R register___U2148 ( .A(register__n4528), .Y(register__n4527) );
  AND2x4_ASAP7_75t_R register___U2149 ( .A(register__n12483), .B(register__n12502), .Y(register__n1963) );
  NAND2x1_ASAP7_75t_R register___U2150 ( .A(register__n516), .B(register__n517), .Y(register__n518) );
  INVxp67_ASAP7_75t_R register___U2151 ( .A(register__n1687), .Y(register__n516) );
  INVxp67_ASAP7_75t_R register___U2152 ( .A(register__net63216), .Y(register__n517) );
  NAND3x1_ASAP7_75t_R register___U2153 ( .A(register__n521), .B(register__n520), .C(register__n522), .Y(register__n519) );
  OA21x2_ASAP7_75t_R register___U2154 ( .A1(register__n112), .A2(register__n2433), .B(register__n2451), .Y(register__n520) );
  OA21x2_ASAP7_75t_R register___U2155 ( .A1(register__net122250), .A2(register__n2430), .B(register__n2449), .Y(register__n521)
         );
  OA21x2_ASAP7_75t_R register___U2156 ( .A1(register__n_cell_124938_net165675), .A2(register__n2431), .B(
        n2450), .Y(register__n522) );
  BUFx12f_ASAP7_75t_R register___U2157 ( .A(register__net143546), .Y(register__net63216) );
  INVx2_ASAP7_75t_R register___U2158 ( .A(register__net96598), .Y(register__n880) );
  INVx2_ASAP7_75t_R register___U2159 ( .A(register__net96598), .Y(register__n2492) );
  HB1xp67_ASAP7_75t_R register___U2160 ( .A(register__C6423_net69274), .Y(register__net128125) );
  BUFx12f_ASAP7_75t_R register___U2161 ( .A(register__net122313), .Y(register__net129787) );
  CKINVDCx20_ASAP7_75t_R register___U2162 ( .A(register__n10285), .Y(register__n523) );
  CKINVDCx5p33_ASAP7_75t_R register___U2163 ( .A(register__n12412), .Y(register__n12401) );
  BUFx6f_ASAP7_75t_R register___U2164 ( .A(register__n3516), .Y(register__n3423) );
  INVx13_ASAP7_75t_R register___U2165 ( .A(register__n2020), .Y(register__n1988) );
  BUFx6f_ASAP7_75t_R register___U2166 ( .A(register__net129017), .Y(register__net102299) );
  BUFx6f_ASAP7_75t_R register___U2167 ( .A(register__n84), .Y(register__net129017) );
  NOR2xp67_ASAP7_75t_R register___U2168 ( .A(register__n12463), .B(register__n4267), .Y(register__n526) );
  NOR2xp33_ASAP7_75t_R register___U2169 ( .A(register__n9055), .B(register__n3708), .Y(register__n527) );
  NOR2xp67_ASAP7_75t_R register___U2170 ( .A(register__n526), .B(register__n527), .Y(register__n12607) );
  HB1xp67_ASAP7_75t_R register___U2171 ( .A(register__n9800), .Y(register__n9055) );
  BUFx6f_ASAP7_75t_R register___U2172 ( .A(register__n11904), .Y(register__n3708) );
  AND2x2_ASAP7_75t_R register___U2173 ( .A(register__n11428), .B(register__n11429), .Y(register__n528) );
  AND4x1_ASAP7_75t_R register___U2174 ( .A(register__n6747), .B(register__n6745), .C(register__n7006), .D(register__n4225), .Y(
        n11429) );
  OAI22xp33_ASAP7_75t_R register___U2175 ( .A1(register__n12401), .A2(register__n460), .B1(register__n10283), .B2(register__n470), 
        .Y(register__n529) );
  CKINVDCx20_ASAP7_75t_R register___U2176 ( .A(register__n10034), .Y(register__n532) );
  INVx2_ASAP7_75t_R register___U2177 ( .A(register__n12353), .Y(register__n12337) );
  INVx1_ASAP7_75t_R register___U2178 ( .A(register__n11100), .Y(register__n533) );
  HB1xp67_ASAP7_75t_R register___U2179 ( .A(register__n11806), .Y(register__n534) );
  HB1xp67_ASAP7_75t_R register___U2180 ( .A(register__n11806), .Y(register__n535) );
  BUFx3_ASAP7_75t_R register___U2181 ( .A(register__n3605), .Y(register__n3261) );
  BUFx6f_ASAP7_75t_R register___U2182 ( .A(register__n12500), .Y(register__n4177) );
  BUFx12f_ASAP7_75t_R register___U2183 ( .A(register__n4920), .Y(register__n3508) );
  BUFx12f_ASAP7_75t_R register___U2184 ( .A(register__n11806), .Y(register__n11804) );
  BUFx6f_ASAP7_75t_R register___U2185 ( .A(register__n3508), .Y(register__n3478) );
  CKINVDCx14_ASAP7_75t_R register___U2186 ( .A(register__n11804), .Y(register__n2220) );
  INVx1_ASAP7_75t_R register___U2187 ( .A(write_data[10]), .Y(register__n861) );
  AND2x2_ASAP7_75t_R register___U2188 ( .A(register__n7675), .B(register__n10974), .Y(register__n536) );
  AND3x1_ASAP7_75t_R register___U2189 ( .A(register__n536), .B(register__n8221), .C(register__n10973), .Y(register__n7024) );
  NAND2xp67_ASAP7_75t_R register___U2190 ( .A(register__n548), .B(register__n538), .Y(register__n545) );
  INVx1_ASAP7_75t_R register___U2191 ( .A(register__n537), .Y(register__n538) );
  INVxp33_ASAP7_75t_R register___U2192 ( .A(register__n627), .Y(register__n539) );
  INVxp33_ASAP7_75t_R register___U2193 ( .A(register__C6423_net61348), .Y(register__n540) );
  INVxp33_ASAP7_75t_R register___U2194 ( .A(register__C6423_net61348), .Y(register__n541) );
  INVxp33_ASAP7_75t_R register___U2195 ( .A(register__n628), .Y(register__n639) );
  INVxp33_ASAP7_75t_R register___U2196 ( .A(register__n630), .Y(register__n635) );
  INVxp33_ASAP7_75t_R register___U2197 ( .A(register__n631), .Y(register__n637) );
  INVxp33_ASAP7_75t_R register___U2198 ( .A(register__n541), .Y(register__n636) );
  INVxp67_ASAP7_75t_R register___U2199 ( .A(register__n631), .Y(register__n642) );
  INVx2_ASAP7_75t_R register___U2200 ( .A(register__n625), .Y(register__n650) );
  INVx2_ASAP7_75t_R register___U2201 ( .A(register__n2022), .Y(register__n625) );
  INVx1_ASAP7_75t_R register___U2202 ( .A(register__n12763), .Y(register__n542) );
  INVxp67_ASAP7_75t_R register___U2203 ( .A(register__n13087), .Y(register__n7077) );
  XNOR2x2_ASAP7_75t_R register___U2204 ( .A(register__n1884), .B(register__n1128), .Y(register__n12518) );
  AOI222xp33_ASAP7_75t_R register___U2205 ( .A1(register__net109611), .A2(register__n9140), .B1(register__net131638), 
        .B2(register__n543), .C1(register__n831), .C2(register__n9217), .Y(register__n11702) );
  INVx3_ASAP7_75t_R register___U2206 ( .A(register__n11710), .Y(register__n7317) );
  HB1xp67_ASAP7_75t_R register___U2207 ( .A(Reg_data[796]), .Y(register__n8095) );
  INVx1_ASAP7_75t_R register___U2208 ( .A(register__n9521), .Y(register__n11664) );
  INVxp33_ASAP7_75t_R register___U2209 ( .A(register__n9521), .Y(register__n1244) );
  INVx2_ASAP7_75t_R register___U2210 ( .A(register__n12493), .Y(register__n1140) );
  INVx3_ASAP7_75t_R register___U2211 ( .A(register__n12493), .Y(register__n1139) );
  INVx1_ASAP7_75t_R register___U2212 ( .A(register__n13270), .Y(register__n4276) );
  BUFx6f_ASAP7_75t_R register___U2213 ( .A(register__n12301), .Y(register__n3358) );
  BUFx6f_ASAP7_75t_R register___U2214 ( .A(register__n12301), .Y(register__n3357) );
  INVx1_ASAP7_75t_R register___U2215 ( .A(register__n12540), .Y(register__n544) );
  OR2x2_ASAP7_75t_R register___U2216 ( .A(register__n2598), .B(register__n2419), .Y(register__n547) );
  OR2x2_ASAP7_75t_R register___U2217 ( .A(register__n1440), .B(register__n2594), .Y(register__n548) );
  INVxp67_ASAP7_75t_R register___U2218 ( .A(register__n3686), .Y(register__n5716) );
  AOI22xp33_ASAP7_75t_R register___U2219 ( .A1(register__n550), .A2(register__net93569), .B1(register__n10173), .B2(
        C6423_net74857), .Y(register__n549) );
  CKINVDCx20_ASAP7_75t_R register___U2220 ( .A(register__n1402), .Y(register__n550) );
  NOR2xp33_ASAP7_75t_R register___U2221 ( .A(register__net127626), .B(register__n6479), .Y(register__n758) );
  OAI22xp5_ASAP7_75t_R register___U2222 ( .A1(register__n53), .A2(register__n7942), .B1(register__net61369), .B2(register__n11965), .Y(read_reg_data_1[1]) );
  INVxp67_ASAP7_75t_R register___U2223 ( .A(register__n845), .Y(register__n12772) );
  OAI22xp33_ASAP7_75t_R register___U2224 ( .A1(register__net63348), .A2(register__n113), .B1(register__n9834), .B2(
        n1541), .Y(register__n551) );
  INVx1_ASAP7_75t_R register___U2225 ( .A(register__n12893), .Y(register__n6188) );
  INVx2_ASAP7_75t_R register___U2226 ( .A(register__n11032), .Y(register__n7606) );
  INVx1_ASAP7_75t_R register___U2227 ( .A(register__n13292), .Y(register__n552) );
  CKINVDCx20_ASAP7_75t_R register___U2228 ( .A(register__n8759), .Y(register__n553) );
  CKINVDCx5p33_ASAP7_75t_R register___U2229 ( .A(register__n3347), .Y(register__n12343) );
  INVx1_ASAP7_75t_R register___U2230 ( .A(register__n5721), .Y(register__n1412) );
  INVxp67_ASAP7_75t_R register___U2231 ( .A(register__n11702), .Y(register__n8322) );
  INVx1_ASAP7_75t_R register___U2232 ( .A(register__n13097), .Y(register__n555) );
  INVx4_ASAP7_75t_R register___U2233 ( .A(n3), .Y(register__n5045) );
  AND2x4_ASAP7_75t_R register___U2234 ( .A(register__n597), .B(register__n7996), .Y(register__C6423_net60462) );
  NAND2xp33_ASAP7_75t_R register___U2235 ( .A(register__n1851), .B(register__n1500), .Y(register__n557) );
  NAND2xp33_ASAP7_75t_R register___U2236 ( .A(register__n556), .B(register__n557), .Y(read_reg_data_1[27]) );
  INVxp67_ASAP7_75t_R register___U2237 ( .A(register__net63028), .Y(register__n1500) );
  HB1xp67_ASAP7_75t_R register___U2238 ( .A(register__n12567), .Y(register__n5976) );
  BUFx6f_ASAP7_75t_R register___U2239 ( .A(register__n11762), .Y(register__n4431) );
  HB1xp67_ASAP7_75t_R register___U2240 ( .A(register__n11553), .Y(register__n4220) );
  HB1xp67_ASAP7_75t_R register___U2241 ( .A(register__n13103), .Y(register__n5792) );
  INVx1_ASAP7_75t_R register___U2242 ( .A(register__n10842), .Y(register__n558) );
  AND2x2_ASAP7_75t_R register___U2243 ( .A(register__n560), .B(register__n2397), .Y(register__n1284) );
  NOR2xp67_ASAP7_75t_R register___U2244 ( .A(register__n559), .B(register__n1285), .Y(register__n560) );
  INVx3_ASAP7_75t_R register___U2245 ( .A(register__net91395), .Y(register__C6422_net59729) );
  NOR2xp33_ASAP7_75t_R register___U2246 ( .A(register__n1335), .B(register__n7697), .Y(register__n1106) );
  HB1xp67_ASAP7_75t_R register___U2247 ( .A(register__n12503), .Y(register__n1904) );
  HB1xp67_ASAP7_75t_R register___U2248 ( .A(register__n3007), .Y(register__n3006) );
  NOR2xp67_ASAP7_75t_R register___U2249 ( .A(register__n1800), .B(register__net113304), .Y(register__n858) );
  INVx1_ASAP7_75t_R register___U2250 ( .A(register__n13368), .Y(register__n562) );
  INVx2_ASAP7_75t_R register___U2251 ( .A(register__n3993), .Y(register__n946) );
  INVx1_ASAP7_75t_R register___U2252 ( .A(register__n4122), .Y(register__n884) );
  INVx1_ASAP7_75t_R register___U2253 ( .A(register__n12779), .Y(register__n563) );
  INVx1_ASAP7_75t_R register___U2254 ( .A(register__n6267), .Y(register__n12421) );
  AOI22xp33_ASAP7_75t_R register___U2255 ( .A1(register__n9351), .A2(register__net110414), .B1(register__n8354), .B2(
        net117889), .Y(register__n1083) );
  AO22x1_ASAP7_75t_R register___U2256 ( .A1(register__n9628), .A2(register__net110414), .B1(register__n10091), .B2(
        n1074), .Y(register__n11256) );
  AO22x1_ASAP7_75t_R register___U2257 ( .A1(register__n9625), .A2(register__net110414), .B1(register__n10088), .B2(
        net117890), .Y(register__n11490) );
  AO22x1_ASAP7_75t_R register___U2258 ( .A1(register__n9632), .A2(register__net110414), .B1(register__n10068), .B2(
        net117890), .Y(register__n11215) );
  AO22x1_ASAP7_75t_R register___U2259 ( .A1(register__n8779), .A2(register__net110414), .B1(register__n9371), .B2(register__n1073), .Y(register__n11722) );
  BUFx6f_ASAP7_75t_R register___U2260 ( .A(register__n554), .Y(register__n3365) );
  INVx2_ASAP7_75t_R register___U2261 ( .A(register__n5990), .Y(register__n9241) );
  INVx3_ASAP7_75t_R register___U2262 ( .A(write_data[21]), .Y(register__n12364) );
  BUFx12f_ASAP7_75t_R register___U2263 ( .A(register__net63016), .Y(register__net141387) );
  INVx1_ASAP7_75t_R register___U2264 ( .A(register__net63034), .Y(register__net63000) );
  INVx2_ASAP7_75t_R register___U2265 ( .A(register__net63034), .Y(register__net63006) );
  INVxp33_ASAP7_75t_R register___U2266 ( .A(register__n11143), .Y(register__n564) );
  BUFx6f_ASAP7_75t_R register___U2267 ( .A(register__n3342), .Y(register__n3316) );
  BUFx6f_ASAP7_75t_R register___U2268 ( .A(register__net63048), .Y(register__net129693) );
  INVx1_ASAP7_75t_R register___U2269 ( .A(register__n5615), .Y(register__n566) );
  BUFx6f_ASAP7_75t_R register___U2270 ( .A(register__n11752), .Y(register__n3339) );
  BUFx6f_ASAP7_75t_R register___U2271 ( .A(register__n11752), .Y(register__n11750) );
  BUFx3_ASAP7_75t_R register___U2272 ( .A(register__n11752), .Y(register__n11747) );
  AOI22xp5_ASAP7_75t_R register___U2273 ( .A1(register__net145522), .A2(register__n567), .B1(register__n568), .B2(register__n569), 
        .Y(register__n12855) );
  CKINVDCx20_ASAP7_75t_R register___U2274 ( .A(register__net90037), .Y(register__n568) );
  INVx13_ASAP7_75t_R register___U2275 ( .A(register__n5838), .Y(register__n569) );
  NAND4xp75_ASAP7_75t_R register___U2276 ( .A(register__n8630), .B(register__n8629), .C(register__n8631), .D(register__n5255), 
        .Y(register__n570) );
  NAND4xp75_ASAP7_75t_R register___U2277 ( .A(register__n7310), .B(register__n3318), .C(register__n7309), .D(register__n7308), 
        .Y(register__n571) );
  INVx2_ASAP7_75t_R register___U2278 ( .A(register__n1966), .Y(register__net150044) );
  INVx1_ASAP7_75t_R register___U2279 ( .A(register__n1967), .Y(register__net150042) );
  INVx1_ASAP7_75t_R register___U2280 ( .A(register__n1966), .Y(register__net150046) );
  INVxp67_ASAP7_75t_R register___U2281 ( .A(register__n1966), .Y(register__n2026) );
  INVx1_ASAP7_75t_R register___U2282 ( .A(register__n1967), .Y(register__net150043) );
  INVxp67_ASAP7_75t_R register___U2283 ( .A(register__net150042), .Y(register__net150051) );
  INVxp67_ASAP7_75t_R register___U2284 ( .A(register__net150046), .Y(register__n1950) );
  INVxp67_ASAP7_75t_R register___U2285 ( .A(register__net150044), .Y(register__net150061) );
  INVxp67_ASAP7_75t_R register___U2286 ( .A(register__net150044), .Y(register__net150059) );
  INVxp67_ASAP7_75t_R register___U2287 ( .A(register__net150044), .Y(register__net150048) );
  HB1xp67_ASAP7_75t_R register___U2288 ( .A(register__n3687), .Y(register__n3686) );
  BUFx6f_ASAP7_75t_R register___U2289 ( .A(register__n11754), .Y(register__n573) );
  BUFx4f_ASAP7_75t_R register___U2290 ( .A(register__n11754), .Y(register__n574) );
  INVx2_ASAP7_75t_R register___U2291 ( .A(register__n4641), .Y(register__n575) );
  INVx2_ASAP7_75t_R register___U2292 ( .A(register__n573), .Y(register__n579) );
  INVx2_ASAP7_75t_R register___U2293 ( .A(register__n573), .Y(register__n580) );
  INVx2_ASAP7_75t_R register___U2294 ( .A(register__n573), .Y(register__n581) );
  INVx2_ASAP7_75t_R register___U2295 ( .A(register__n573), .Y(register__n582) );
  INVx2_ASAP7_75t_R register___U2296 ( .A(register__n573), .Y(register__n583) );
  INVx2_ASAP7_75t_R register___U2297 ( .A(register__n573), .Y(register__n584) );
  INVx2_ASAP7_75t_R register___U2298 ( .A(register__n574), .Y(register__n585) );
  INVx2_ASAP7_75t_R register___U2299 ( .A(register__n574), .Y(register__n586) );
  INVx1_ASAP7_75t_R register___U2300 ( .A(register__n574), .Y(register__n587) );
  INVx1_ASAP7_75t_R register___U2301 ( .A(register__n574), .Y(register__n588) );
  INVx1_ASAP7_75t_R register___U2302 ( .A(register__n574), .Y(register__n589) );
  INVx1_ASAP7_75t_R register___U2303 ( .A(register__n574), .Y(register__n590) );
  NAND2xp67_ASAP7_75t_R register___U2304 ( .A(register__net129787), .B(register__net89741), .Y(register__n2450) );
  INVxp67_ASAP7_75t_R register___U2305 ( .A(register__n4142), .Y(register__n9401) );
  INVx1_ASAP7_75t_R register___U2306 ( .A(register__n12971), .Y(register__n591) );
  INVx1_ASAP7_75t_R register___U2307 ( .A(register__n11409), .Y(register__n592) );
  HB1xp67_ASAP7_75t_R register___U2308 ( .A(register__n3543), .Y(register__n4636) );
  CKINVDCx10_ASAP7_75t_R register___U2309 ( .A(register__n12418), .Y(register__n12405) );
  BUFx12f_ASAP7_75t_R register___U2310 ( .A(register__n12419), .Y(register__n12418) );
  BUFx3_ASAP7_75t_R register___U2311 ( .A(register__net99590), .Y(register__net124704) );
  BUFx3_ASAP7_75t_R register___U2312 ( .A(register__n783), .Y(register__net99590) );
  INVxp33_ASAP7_75t_R register___U2313 ( .A(register__net122579), .Y(register__n914) );
  HB1xp67_ASAP7_75t_R register___U2314 ( .A(register__n3782), .Y(register__n3781) );
  AND2x4_ASAP7_75t_R register___U2315 ( .A(register__n385), .B(register__n7684), .Y(register__n12497) );
  INVxp67_ASAP7_75t_R register___U2316 ( .A(register__n12498), .Y(register__n2804) );
  INVx4_ASAP7_75t_R register___U2317 ( .A(register__net63026), .Y(register__net62990) );
  HB1xp67_ASAP7_75t_R register___U2318 ( .A(register__n13387), .Y(register__n4008) );
  BUFx3_ASAP7_75t_R register___U2319 ( .A(register__n3606), .Y(register__n8335) );
  INVxp33_ASAP7_75t_R register___U2320 ( .A(register__net122579), .Y(register__n913) );
  INVxp67_ASAP7_75t_R register___U2321 ( .A(register__n12730), .Y(register__n5719) );
  INVx1_ASAP7_75t_R register___U2322 ( .A(register__n2134), .Y(register__n1745) );
  NOR2xp67_ASAP7_75t_R register___U2323 ( .A(register__n223), .B(register__n1159), .Y(register__n7021) );
  NAND2xp67_ASAP7_75t_R register___U2324 ( .A(register__n7593), .B(register__n2212), .Y(register__n1159) );
  OAI22xp5_ASAP7_75t_R register___U2325 ( .A1(register__net66302), .A2(register__n8641), .B1(register__n4377), .B2(
        n1687), .Y(read_reg_data_2[0]) );
  BUFx6f_ASAP7_75t_R register___U2326 ( .A(register__n11981), .Y(register__n9407) );
  AND4x1_ASAP7_75t_R register___U2327 ( .A(register__n5534), .B(register__n5532), .C(register__n6546), .D(register__n3863), .Y(
        n10995) );
  HB1xp67_ASAP7_75t_R register___U2328 ( .A(register__n12745), .Y(register__n3578) );
  INVx1_ASAP7_75t_R register___U2329 ( .A(register__n12595), .Y(register__n595) );
  HB1xp67_ASAP7_75t_R register___U2330 ( .A(register__n12906), .Y(register__n3007) );
  BUFx6f_ASAP7_75t_R register___U2331 ( .A(register__n12248), .Y(register__n4967) );
  BUFx3_ASAP7_75t_R register___U2332 ( .A(register__n12248), .Y(register__n4839) );
  BUFx6f_ASAP7_75t_R register___U2333 ( .A(register__n3648), .Y(register__n12269) );
  INVxp33_ASAP7_75t_R register___U2334 ( .A(WB_rd[4]), .Y(register__n596) );
  INVxp67_ASAP7_75t_R register___U2335 ( .A(WB_rd[4]), .Y(register__n666) );
  OAI22xp33_ASAP7_75t_R register___U2336 ( .A1(register__n1883), .A2(register__n_cell_125487_net184714), .B1(
        n664), .B2(register__net109643), .Y(register__n10602) );
  INVx2_ASAP7_75t_R register___U2337 ( .A(rs2[1]), .Y(register__n11709) );
  OAI22xp5_ASAP7_75t_R register___U2338 ( .A1(register__net66308), .A2(register__n9154), .B1(register__n12178), .B2(
        n1687), .Y(read_reg_data_2[14]) );
  INVx2_ASAP7_75t_R register___U2339 ( .A(register__n716), .Y(register__n717) );
  AOI22x1_ASAP7_75t_R register___U2340 ( .A1(register__net62706), .A2(register__n598), .B1(register__n599), .B2(register__n600), 
        .Y(register__n12553) );
  CKINVDCx20_ASAP7_75t_R register___U2341 ( .A(register__n9861), .Y(register__n599) );
  CKINVDCx5p33_ASAP7_75t_R register___U2342 ( .A(register__net62706), .Y(register__net62676) );
  BUFx2_ASAP7_75t_R register___U2343 ( .A(register__n3300), .Y(register__n12383) );
  INVx1_ASAP7_75t_R register___U2344 ( .A(register__n12383), .Y(register__n12369) );
  AO22x1_ASAP7_75t_R register___U2345 ( .A1(register__n9646), .A2(register__n3), .B1(register__n9973), .B2(register__n233), .Y(
        n10882) );
  HB1xp67_ASAP7_75t_R register___U2346 ( .A(register__n4141), .Y(register__n4140) );
  HB1xp67_ASAP7_75t_R register___U2347 ( .A(register__n4518), .Y(register__n4517) );
  BUFx6f_ASAP7_75t_R register___U2348 ( .A(register__n12141), .Y(register__n4634) );
  INVx1_ASAP7_75t_R register___U2349 ( .A(register__n12868), .Y(register__n602) );
  INVxp33_ASAP7_75t_R register___U2350 ( .A(register__net114452), .Y(register__n2375) );
  INVxp33_ASAP7_75t_R register___U2351 ( .A(register__n4157), .Y(register__n4278) );
  BUFx2_ASAP7_75t_R register___U2352 ( .A(register__n2803), .Y(register__n2812) );
  HB1xp67_ASAP7_75t_R register___U2353 ( .A(register__n13319), .Y(register__n4528) );
  AND2x4_ASAP7_75t_R register___U2354 ( .A(register__n1963), .B(register__n12485), .Y(register__n12494) );
  INVx1_ASAP7_75t_R register___U2355 ( .A(register__n12957), .Y(register__n604) );
  AOI21xp33_ASAP7_75t_R register___U2356 ( .A1(register__net94399), .A2(register__net89277), .B(register__n2488), .Y(
        n2509) );
  AO22x1_ASAP7_75t_R register___U2357 ( .A1(register__net90937), .A2(register__net125170), .B1(register__net90081), 
        .B2(register__n436), .Y(register__n11286) );
  AO22x1_ASAP7_75t_R register___U2358 ( .A1(register__n9746), .A2(register__net125170), .B1(register__n8455), .B2(register__n515), 
        .Y(register__n11395) );
  AO22x1_ASAP7_75t_R register___U2359 ( .A1(register__n9909), .A2(register__net125170), .B1(register__n6930), .B2(
        C6423_net68914), .Y(register__n11689) );
  AO22x1_ASAP7_75t_R register___U2360 ( .A1(register__n7391), .A2(register__net125170), .B1(register__n4960), .B2(register__n515), 
        .Y(register__n11711) );
  AO22x1_ASAP7_75t_R register___U2361 ( .A1(register__n6285), .A2(register__net125170), .B1(register__n4758), .B2(register__n515), 
        .Y(register__n11569) );
  AO22x1_ASAP7_75t_R register___U2362 ( .A1(register__n8753), .A2(register__net125170), .B1(register__n10229), .B2(register__n515), .Y(register__n11375) );
  INVx1_ASAP7_75t_R register___U2363 ( .A(register__n12958), .Y(register__n607) );
  INVx4_ASAP7_75t_R register___U2364 ( .A(n4), .Y(register__n12079) );
  INVx1_ASAP7_75t_R register___U2365 ( .A(register__n12733), .Y(register__n609) );
  BUFx6f_ASAP7_75t_R register___U2366 ( .A(register__n11751), .Y(register__n2886) );
  BUFx12f_ASAP7_75t_R register___U2367 ( .A(register__n2882), .Y(register__n11751) );
  AO22x1_ASAP7_75t_R register___U2368 ( .A1(register__n9335), .A2(register__net109204), .B1(register__n9355), .B2(
        net129911), .Y(register__n10834) );
  AO22x1_ASAP7_75t_R register___U2369 ( .A1(register__n8193), .A2(register__C6422_net60415), .B1(register__n10233), 
        .B2(register__net88727), .Y(register__n10750) );
  AO22x1_ASAP7_75t_R register___U2370 ( .A1(register__n8104), .A2(register__C6422_net60415), .B1(register__n6112), .B2(
        net88727), .Y(register__n10774) );
  AO22x1_ASAP7_75t_R register___U2371 ( .A1(register__net90669), .A2(register__C6422_net60415), .B1(register__net89593), 
        .B2(register__net88727), .Y(register__n10728) );
  AO22x1_ASAP7_75t_R register___U2372 ( .A1(register__n9674), .A2(register__C6422_net60415), .B1(register__n9921), .B2(
        net88727), .Y(register__n10878) );
  NOR2xp67_ASAP7_75t_R register___U2373 ( .A(register__n12175), .B(register__n179), .Y(register__n2082) );
  NOR2xp67_ASAP7_75t_R register___U2374 ( .A(register__n2082), .B(register__n2083), .Y(register__n12678) );
  AND2x2_ASAP7_75t_R register___U2375 ( .A(register__n11098), .B(register__n11097), .Y(register__n611) );
  AND3x1_ASAP7_75t_R register___U2376 ( .A(register__n611), .B(register__n1271), .C(register__n8261), .Y(register__n8642) );
  HB1xp67_ASAP7_75t_R register___U2377 ( .A(register__n443), .Y(register__n612) );
  OAI22xp33_ASAP7_75t_R register___U2378 ( .A1(register__n12422), .A2(register__n11868), .B1(register__n8548), .B2(
        n11752), .Y(register__n613) );
  BUFx12f_ASAP7_75t_R register___U2379 ( .A(register__n8564), .Y(register__n8561) );
  INVx2_ASAP7_75t_R register___U2380 ( .A(register__n3524), .Y(register__n1050) );
  BUFx6f_ASAP7_75t_R register___U2381 ( .A(register__n6752), .Y(register__n3524) );
  INVx2_ASAP7_75t_R register___U2382 ( .A(register__n3522), .Y(register__n6752) );
  INVxp67_ASAP7_75t_R register___U2383 ( .A(register__n12214), .Y(register__n12194) );
  INVx1_ASAP7_75t_R register___U2384 ( .A(register__n12220), .Y(register__n12203) );
  INVx1_ASAP7_75t_R register___U2385 ( .A(register__n12626), .Y(register__n614) );
  NOR2xp33_ASAP7_75t_R register___U2386 ( .A(register__net98849), .B(register__n1161), .Y(register__n616) );
  INVxp67_ASAP7_75t_R register___U2387 ( .A(register__n13300), .Y(register__n617) );
  BUFx12f_ASAP7_75t_R register___U2388 ( .A(register__net98851), .Y(register__net98849) );
  INVx1_ASAP7_75t_R register___U2389 ( .A(register__n12689), .Y(register__n618) );
  INVxp67_ASAP7_75t_R register___U2390 ( .A(register__n12747), .Y(register__n8582) );
  HB1xp67_ASAP7_75t_R register___U2391 ( .A(register__n5579), .Y(register__n5578) );
  INVx6_ASAP7_75t_R register___U2392 ( .A(register__n6462), .Y(register__n1641) );
  BUFx12f_ASAP7_75t_R register___U2393 ( .A(register__net129692), .Y(register__net129690) );
  BUFx12f_ASAP7_75t_R register___U2394 ( .A(register__net63048), .Y(register__net129692) );
  BUFx3_ASAP7_75t_R register___U2395 ( .A(register__n4867), .Y(register__n4196) );
  BUFx3_ASAP7_75t_R register___U2396 ( .A(register__n4867), .Y(register__n4194) );
  BUFx6f_ASAP7_75t_R register___U2397 ( .A(register__n4867), .Y(register__n4193) );
  BUFx12f_ASAP7_75t_R register___U2398 ( .A(register__n12050), .Y(register__n4867) );
  INVx1_ASAP7_75t_R register___U2399 ( .A(register__n12851), .Y(register__n619) );
  INVx1_ASAP7_75t_R register___U2400 ( .A(register__n3832), .Y(register__n11810) );
  BUFx12f_ASAP7_75t_R register___U2401 ( .A(register__n3705), .Y(register__n3507) );
  NOR2xp33_ASAP7_75t_R register___U2402 ( .A(register__n2002), .B(register__n5729), .Y(register__n620) );
  NOR3xp33_ASAP7_75t_R register___U2403 ( .A(register__n620), .B(register__n621), .C(register__n622), .Y(register__n10526) );
  AND2x2_ASAP7_75t_R register___U2404 ( .A(register__n10524), .B(register__n10523), .Y(register__n623) );
  AND3x1_ASAP7_75t_R register___U2405 ( .A(register__n623), .B(register__n8565), .C(register__n8302), .Y(register__n9180) );
  HB1xp67_ASAP7_75t_R register___U2406 ( .A(register__n10532), .Y(register__n5729) );
  BUFx3_ASAP7_75t_R register___U2407 ( .A(register__n10533), .Y(register__n7580) );
  HB1xp67_ASAP7_75t_R register___U2408 ( .A(register__n10534), .Y(register__n6469) );
  BUFx2_ASAP7_75t_R register___U2409 ( .A(register__n10522), .Y(register__n8565) );
  INVx1_ASAP7_75t_R register___U2410 ( .A(register__n5125), .Y(register__n8302) );
  BUFx6f_ASAP7_75t_R register___U2411 ( .A(register__n12164), .Y(register__n3256) );
  BUFx6f_ASAP7_75t_R register___U2412 ( .A(register__n3256), .Y(register__n3254) );
  INVx1_ASAP7_75t_R register___U2413 ( .A(register__n12636), .Y(register__n624) );
  INVxp67_ASAP7_75t_R register___U2414 ( .A(register__n4298), .Y(register__n7617) );
  INVxp67_ASAP7_75t_R register___U2415 ( .A(register__n3742), .Y(register__n5712) );
  NAND2xp5_ASAP7_75t_R register___U2416 ( .A(register__net146144), .B(register__net96895), .Y(register__n2353) );
  HB1xp67_ASAP7_75t_R register___U2417 ( .A(register__n4106), .Y(register__n4105) );
  INVxp33_ASAP7_75t_R register___U2418 ( .A(register__C6423_net61348), .Y(register__n626) );
  INVxp67_ASAP7_75t_R register___U2419 ( .A(register__C6423_net61348), .Y(register__n627) );
  INVxp67_ASAP7_75t_R register___U2420 ( .A(register__C6423_net61348), .Y(register__n628) );
  INVxp33_ASAP7_75t_R register___U2421 ( .A(register__C6423_net61348), .Y(register__n629) );
  INVxp33_ASAP7_75t_R register___U2422 ( .A(register__C6423_net61348), .Y(register__n630) );
  INVxp33_ASAP7_75t_R register___U2423 ( .A(register__n627), .Y(register__n632) );
  INVxp33_ASAP7_75t_R register___U2424 ( .A(register__n629), .Y(register__n633) );
  INVxp33_ASAP7_75t_R register___U2425 ( .A(register__n626), .Y(register__n634) );
  INVxp33_ASAP7_75t_R register___U2426 ( .A(register__n628), .Y(register__n638) );
  INVxp67_ASAP7_75t_R register___U2427 ( .A(register__n628), .Y(register__n640) );
  INVxp33_ASAP7_75t_R register___U2428 ( .A(register__n630), .Y(register__n641) );
  INVxp33_ASAP7_75t_R register___U2429 ( .A(register__n540), .Y(register__n643) );
  INVxp33_ASAP7_75t_R register___U2430 ( .A(register__n541), .Y(register__n644) );
  INVxp33_ASAP7_75t_R register___U2431 ( .A(register__n630), .Y(register__n645) );
  INVxp33_ASAP7_75t_R register___U2432 ( .A(register__n627), .Y(register__n646) );
  INVxp33_ASAP7_75t_R register___U2433 ( .A(register__n629), .Y(register__n647) );
  INVxp33_ASAP7_75t_R register___U2434 ( .A(register__n626), .Y(register__n648) );
  INVxp33_ASAP7_75t_R register___U2435 ( .A(register__n540), .Y(register__n649) );
  BUFx2_ASAP7_75t_R register___U2436 ( .A(register__C6423_net61348), .Y(register__n2022) );
  BUFx6f_ASAP7_75t_R register___U2437 ( .A(register__n11813), .Y(register__n3308) );
  BUFx6f_ASAP7_75t_R register___U2438 ( .A(register__net147144), .Y(register__net125383) );
  INVx1_ASAP7_75t_R register___U2439 ( .A(register__n13281), .Y(register__n5937) );
  BUFx12f_ASAP7_75t_R register___U2440 ( .A(register__n3909), .Y(register__n3276) );
  HB1xp67_ASAP7_75t_R register___U2441 ( .A(register__n12949), .Y(register__n5754) );
  INVx2_ASAP7_75t_R register___U2442 ( .A(register__n11236), .Y(register__n8233) );
  INVx2_ASAP7_75t_R register___U2443 ( .A(register__n1081), .Y(register__n1082) );
  AND2x2_ASAP7_75t_R register___U2444 ( .A(register__n12483), .B(register__n12502), .Y(register__n12492) );
  INVxp67_ASAP7_75t_R register___U2445 ( .A(register__n11813), .Y(register__n1100) );
  INVxp67_ASAP7_75t_R register___U2446 ( .A(register__n11813), .Y(register__n1633) );
  AND3x1_ASAP7_75t_R register___U2447 ( .A(register__n1477), .B(register__n2903), .C(register__n1222), .Y(register__n8250) );
  INVx2_ASAP7_75t_R register___U2448 ( .A(register__n3343), .Y(register__n708) );
  BUFx6f_ASAP7_75t_R register___U2449 ( .A(register__net62690), .Y(register__net144153) );
  INVx2_ASAP7_75t_R register___U2450 ( .A(register__net62690), .Y(register__net62658) );
  BUFx6f_ASAP7_75t_R register___U2451 ( .A(register__net141449), .Y(register__net62690) );
  BUFx6f_ASAP7_75t_R register___U2452 ( .A(register__net144153), .Y(register__net121463) );
  INVxp67_ASAP7_75t_R register___U2453 ( .A(register__n12379), .Y(register__n3467) );
  INVx1_ASAP7_75t_R register___U2454 ( .A(register__n12379), .Y(register__n12365) );
  INVxp67_ASAP7_75t_R register___U2455 ( .A(register__n12387), .Y(register__n12372) );
  INVx3_ASAP7_75t_R register___U2456 ( .A(register__C6423_net68920), .Y(register__n2419) );
  BUFx4f_ASAP7_75t_R register___U2457 ( .A(register__net128121), .Y(register__C6423_net68920) );
  INVx1_ASAP7_75t_R register___U2458 ( .A(register__n12768), .Y(register__n2250) );
  NOR2x1p5_ASAP7_75t_R register___U2459 ( .A(register__n2782), .B(register__n2783), .Y(register__n12768) );
  NOR2x2_ASAP7_75t_R register___U2460 ( .A(register__n12060), .B(register__n115), .Y(register__n2782) );
  HB1xp67_ASAP7_75t_R register___U2461 ( .A(Reg_data[476]), .Y(register__n9065) );
  INVx1_ASAP7_75t_R register___U2462 ( .A(register__n2938), .Y(register__n1375) );
  BUFx6f_ASAP7_75t_R register___U2463 ( .A(register__n11760), .Y(register__n7336) );
  BUFx12f_ASAP7_75t_R register___U2464 ( .A(register__n5531), .Y(register__n11760) );
  NAND3xp33_ASAP7_75t_R register___U2465 ( .A(register__n406), .B(register__n5441), .C(register__n11721), .Y(register__n652) );
  HB1xp67_ASAP7_75t_R register___U2466 ( .A(register__n4143), .Y(register__n4142) );
  BUFx12f_ASAP7_75t_R register___U2467 ( .A(register__net143813), .Y(register__net143812) );
  HB1xp67_ASAP7_75t_R register___U2468 ( .A(register__n3246), .Y(register__n3245) );
  OAI22xp33_ASAP7_75t_R register___U2469 ( .A1(register__net62652), .A2(register__n1049), .B1(register__n7843), .B2(
        n3276), .Y(register__n654) );
  INVxp67_ASAP7_75t_R register___U2470 ( .A(register__n3028), .Y(register__n3942) );
  HB1xp67_ASAP7_75t_R register___U2471 ( .A(register__n3029), .Y(register__n3028) );
  NOR3x1_ASAP7_75t_R register___U2472 ( .A(register__n21), .B(register__n5606), .C(register__n1854), .Y(register__n11034) );
  AO22x1_ASAP7_75t_R register___U2473 ( .A1(register__n9706), .A2(register__net129017), .B1(register__n10036), .B2(register__n422), .Y(register__n11534) );
  AO22x1_ASAP7_75t_R register___U2474 ( .A1(register__n8910), .A2(register__net129017), .B1(register__n10048), .B2(register__n422), .Y(register__n11213) );
  AO22x1_ASAP7_75t_R register___U2475 ( .A1(register__net95451), .A2(register__net129017), .B1(register__net89817), 
        .B2(register__n422), .Y(register__n11291) );
  HB1xp67_ASAP7_75t_R register___U2476 ( .A(register__n13041), .Y(register__n5088) );
  BUFx3_ASAP7_75t_R register___U2477 ( .A(register__net129692), .Y(register__net63036) );
  AOI22x1_ASAP7_75t_R register___U2478 ( .A1(register__n12000), .A2(register__n656), .B1(register__n657), .B2(register__n658), 
        .Y(register__n13386) );
  CKINVDCx20_ASAP7_75t_R register___U2479 ( .A(register__n11730), .Y(register__n656) );
  CKINVDCx20_ASAP7_75t_R register___U2480 ( .A(register__n10359), .Y(register__n657) );
  CKINVDCx20_ASAP7_75t_R register___U2481 ( .A(register__n1164), .Y(register__n658) );
  INVx2_ASAP7_75t_R register___U2482 ( .A(register__n12000), .Y(register__n11983) );
  HB1xp67_ASAP7_75t_R register___U2483 ( .A(register__n12775), .Y(register__n4500) );
  NAND2xp67_ASAP7_75t_R register___U2484 ( .A(register__n641), .B(register__net88496), .Y(register__n2522) );
  AO22x1_ASAP7_75t_R register___U2485 ( .A1(register__n9654), .A2(register__net109849), .B1(register__n9981), .B2(register__n646), 
        .Y(register__n11218) );
  AND2x2_ASAP7_75t_R register___U2486 ( .A(rs2[0]), .B(register__n11709), .Y(register__n2744) );
  INVx1_ASAP7_75t_R register___U2487 ( .A(register__n12948), .Y(register__n659) );
  HB1xp67_ASAP7_75t_R register___U2488 ( .A(register__n2881), .Y(register__n3275) );
  INVxp67_ASAP7_75t_R register___U2489 ( .A(register__n6250), .Y(register__n9184) );
  HB1xp67_ASAP7_75t_R register___U2490 ( .A(register__n12418), .Y(register__n5350) );
  OAI22xp33_ASAP7_75t_R register___U2491 ( .A1(register__n12342), .A2(register__n893), .B1(register__n9660), .B2(register__n899), 
        .Y(register__n661) );
  INVx1_ASAP7_75t_R register___U2492 ( .A(register__n13019), .Y(register__n662) );
  BUFx6f_ASAP7_75t_R register___U2493 ( .A(register__n3265), .Y(register__n3283) );
  INVx6_ASAP7_75t_R register___U2494 ( .A(register__n12212), .Y(register__n12197) );
  BUFx12f_ASAP7_75t_R register___U2495 ( .A(register__n3364), .Y(register__n12212) );
  BUFx6f_ASAP7_75t_R register___U2496 ( .A(register__n9407), .Y(register__n11969) );
  HB1xp67_ASAP7_75t_R register___U2497 ( .A(register__n10673), .Y(register__n4106) );
  BUFx3_ASAP7_75t_R register___U2498 ( .A(register__n3268), .Y(register__n11812) );
  INVxp67_ASAP7_75t_R register___U2499 ( .A(register__n3268), .Y(register__n1783) );
  HB1xp67_ASAP7_75t_R register___U2500 ( .A(register__n4406), .Y(register__n4405) );
  BUFx3_ASAP7_75t_R register___U2501 ( .A(register__n3023), .Y(register__n3004) );
  BUFx6f_ASAP7_75t_R register___U2502 ( .A(register__n12277), .Y(register__n3070) );
  AND2x4_ASAP7_75t_R register___U2503 ( .A(register__n389), .B(register__n740), .Y(register__C6423_net60464) );
  BUFx6f_ASAP7_75t_R register___U2504 ( .A(register__n3628), .Y(register__n12135) );
  CKINVDCx20_ASAP7_75t_R register___U2505 ( .A(register__n9547), .Y(register__n663) );
  HB1xp67_ASAP7_75t_R register___U2506 ( .A(register__n4396), .Y(register__n4395) );
  CKINVDCx5p33_ASAP7_75t_R register___U2507 ( .A(register__n12044), .Y(register__n12028) );
  BUFx12f_ASAP7_75t_R register___U2508 ( .A(register__n4728), .Y(register__n12412) );
  HB1xp67_ASAP7_75t_R register___U2509 ( .A(register__n4299), .Y(register__n4298) );
  INVxp67_ASAP7_75t_R register___U2510 ( .A(register__n2987), .Y(register__n4985) );
  HB1xp67_ASAP7_75t_R register___U2511 ( .A(register__n2988), .Y(register__n2987) );
  HB1xp67_ASAP7_75t_R register___U2512 ( .A(register__n6251), .Y(register__n6250) );
  INVxp67_ASAP7_75t_R register___U2513 ( .A(register__n3655), .Y(register__n6732) );
  BUFx6f_ASAP7_75t_R register___U2514 ( .A(register__n12364), .Y(register__n5349) );
  HB1xp67_ASAP7_75t_R register___U2515 ( .A(register__n12556), .Y(register__n4602) );
  BUFx6f_ASAP7_75t_R register___U2516 ( .A(register__n4290), .Y(register__n7906) );
  BUFx12f_ASAP7_75t_R register___U2517 ( .A(register__n12079), .Y(register__n12078) );
  NOR2x1_ASAP7_75t_R register___U2518 ( .A(register__n2275), .B(register__n2276), .Y(register__n1081) );
  NAND4xp75_ASAP7_75t_R register___U2519 ( .A(register__n7317), .B(register__n7315), .C(register__n8265), .D(register__n4256), 
        .Y(register__n2276) );
  INVxp67_ASAP7_75t_R register___U2520 ( .A(register__n1490), .Y(register__n12936) );
  AO22x1_ASAP7_75t_R register___U2521 ( .A1(register__n12164), .A2(register__n474), .B1(register__n1491), .B2(register__n461), 
        .Y(register__n1490) );
  BUFx2_ASAP7_75t_R register___U2522 ( .A(register__n667), .Y(register__net141508) );
  NAND3x1_ASAP7_75t_R register___U2523 ( .A(register__n11451), .B(register__n11452), .C(register__n11453), .Y(register__n11450)
         );
  INVxp67_ASAP7_75t_R register___U2524 ( .A(register__n2951), .Y(register__n4645) );
  BUFx4f_ASAP7_75t_R register___U2525 ( .A(register__n3570), .Y(register__n3568) );
  INVx3_ASAP7_75t_R register___U2526 ( .A(register__n12477), .Y(register__n12464) );
  HB1xp67_ASAP7_75t_R register___U2527 ( .A(register__n12920), .Y(register__n5784) );
  BUFx3_ASAP7_75t_R register___U2528 ( .A(register__n3918), .Y(register__n3511) );
  BUFx12f_ASAP7_75t_R register___U2529 ( .A(register__n11763), .Y(register__n5173) );
  INVxp67_ASAP7_75t_R register___U2530 ( .A(register__n1847), .Y(register__n668) );
  INVxp67_ASAP7_75t_R register___U2531 ( .A(register__n1845), .Y(register__n669) );
  INVxp67_ASAP7_75t_R register___U2532 ( .A(register__n1846), .Y(register__n670) );
  INVxp67_ASAP7_75t_R register___U2533 ( .A(register__n1844), .Y(register__n671) );
  INVxp67_ASAP7_75t_R register___U2534 ( .A(register__n1843), .Y(register__n672) );
  INVxp67_ASAP7_75t_R register___U2535 ( .A(register__n1849), .Y(register__n673) );
  INVxp33_ASAP7_75t_R register___U2536 ( .A(register__n11740), .Y(register__n674) );
  INVxp67_ASAP7_75t_R register___U2537 ( .A(register__n811), .Y(register__n675) );
  INVxp67_ASAP7_75t_R register___U2538 ( .A(register__n808), .Y(register__n676) );
  INVxp67_ASAP7_75t_R register___U2539 ( .A(register__n807), .Y(register__n677) );
  INVxp33_ASAP7_75t_R register___U2540 ( .A(register__n812), .Y(register__n678) );
  INVxp67_ASAP7_75t_R register___U2541 ( .A(register__n810), .Y(register__n679) );
  INVx2_ASAP7_75t_R register___U2542 ( .A(register__n4475), .Y(register__n680) );
  INVx1_ASAP7_75t_R register___U2543 ( .A(register__n4476), .Y(register__n681) );
  INVx1_ASAP7_75t_R register___U2544 ( .A(register__n1901), .Y(register__n682) );
  INVx1_ASAP7_75t_R register___U2545 ( .A(register__n11739), .Y(register__n683) );
  INVx1_ASAP7_75t_R register___U2546 ( .A(register__n2945), .Y(register__n684) );
  INVx2_ASAP7_75t_R register___U2547 ( .A(register__n11738), .Y(register__n685) );
  INVx1_ASAP7_75t_R register___U2548 ( .A(register__n11853), .Y(register__n686) );
  INVx1_ASAP7_75t_R register___U2549 ( .A(register__n11854), .Y(register__n687) );
  INVx6_ASAP7_75t_R register___U2550 ( .A(register__n3075), .Y(register__n688) );
  INVx6_ASAP7_75t_R register___U2551 ( .A(register__n11737), .Y(register__n689) );
  INVx1_ASAP7_75t_R register___U2552 ( .A(register__n11855), .Y(register__n690) );
  INVx1_ASAP7_75t_R register___U2553 ( .A(register__n11857), .Y(register__n691) );
  INVx1_ASAP7_75t_R register___U2554 ( .A(register__n11856), .Y(register__n692) );
  INVx2_ASAP7_75t_R register___U2555 ( .A(register__n3074), .Y(register__n693) );
  INVx1_ASAP7_75t_R register___U2556 ( .A(register__n814), .Y(register__n694) );
  INVx1_ASAP7_75t_R register___U2557 ( .A(register__n813), .Y(register__n695) );
  INVx1_ASAP7_75t_R register___U2558 ( .A(register__n816), .Y(register__n696) );
  INVx1_ASAP7_75t_R register___U2559 ( .A(register__n815), .Y(register__n697) );
  INVx2_ASAP7_75t_R register___U2560 ( .A(register__n4851), .Y(register__n699) );
  INVx2_ASAP7_75t_R register___U2561 ( .A(register__n4851), .Y(register__n700) );
  INVx1_ASAP7_75t_R register___U2562 ( .A(register__n4851), .Y(register__n702) );
  BUFx4f_ASAP7_75t_R register___U2563 ( .A(register__n4851), .Y(register__n11858) );
  BUFx6f_ASAP7_75t_R register___U2564 ( .A(register__n11858), .Y(register__n2163) );
  BUFx3_ASAP7_75t_R register___U2565 ( .A(register__n4851), .Y(register__n806) );
  INVx6_ASAP7_75t_R register___U2566 ( .A(register__n11858), .Y(register__n11740) );
  BUFx12f_ASAP7_75t_R register___U2567 ( .A(register__n11740), .Y(register__n4476) );
  BUFx12f_ASAP7_75t_R register___U2568 ( .A(register__n4476), .Y(register__n2945) );
  INVx1_ASAP7_75t_R register___U2569 ( .A(register__n3868), .Y(register__n11855) );
  BUFx4f_ASAP7_75t_R register___U2570 ( .A(register__n11739), .Y(register__n3074) );
  INVx1_ASAP7_75t_R register___U2571 ( .A(register__n806), .Y(register__n814) );
  INVx1_ASAP7_75t_R register___U2572 ( .A(register__n806), .Y(register__n813) );
  INVx1_ASAP7_75t_R register___U2573 ( .A(register__n806), .Y(register__n816) );
  INVx1_ASAP7_75t_R register___U2574 ( .A(register__n806), .Y(register__n815) );
  INVx2_ASAP7_75t_R register___U2575 ( .A(register__n11827), .Y(register__n2286) );
  BUFx6f_ASAP7_75t_R register___U2576 ( .A(register__n12141), .Y(register__n3543) );
  HB1xp67_ASAP7_75t_R register___U2577 ( .A(register__n12989), .Y(register__n4157) );
  HB1xp67_ASAP7_75t_R register___U2578 ( .A(register__n3660), .Y(register__n3659) );
  AND4x1_ASAP7_75t_R register___U2579 ( .A(register__n1325), .B(register__n7054), .C(register__n7055), .D(register__n5394), .Y(
        n11321) );
  BUFx3_ASAP7_75t_R register___U2580 ( .A(register__net63054), .Y(register__net136188) );
  BUFx6f_ASAP7_75t_R register___U2581 ( .A(register__net64864), .Y(register__net64900) );
  AO22x1_ASAP7_75t_R register___U2582 ( .A1(register__n9682), .A2(register__C6422_net60422), .B1(register__n9953), .B2(
        net123857), .Y(register__n10966) );
  BUFx6f_ASAP7_75t_R register___U2583 ( .A(register__n11947), .Y(register__n11946) );
  NOR2xp33_ASAP7_75t_R register___U2584 ( .A(register__n786), .B(register__n785), .Y(register__n703) );
  NOR2xp33_ASAP7_75t_R register___U2585 ( .A(register__n787), .B(register__n704), .Y(register__n4950) );
  INVxp33_ASAP7_75t_R register___U2586 ( .A(register__n703), .Y(register__n704) );
  NOR2xp33_ASAP7_75t_R register___U2587 ( .A(register__net112578), .B(register__n6473), .Y(register__n787) );
  NOR2x1_ASAP7_75t_R register___U2588 ( .A(register__n1047), .B(register__n1048), .Y(register__n7888) );
  BUFx4f_ASAP7_75t_R register___U2589 ( .A(register__n1762), .Y(register__n7697) );
  BUFx3_ASAP7_75t_R register___U2590 ( .A(register__n5501), .Y(register__n8358) );
  INVxp67_ASAP7_75t_R register___U2591 ( .A(register__n3394), .Y(register__n4384) );
  HB1xp67_ASAP7_75t_R register___U2592 ( .A(register__n3395), .Y(register__n3394) );
  INVxp67_ASAP7_75t_R register___U2593 ( .A(register__n10877), .Y(register__n8571) );
  BUFx12f_ASAP7_75t_R register___U2594 ( .A(register__n3268), .Y(register__n11813) );
  OAI22xp5_ASAP7_75t_R register___U2595 ( .A1(register__n54), .A2(register__n3720), .B1(register__net61369), .B2(register__n12164), .Y(read_reg_data_1[13]) );
  INVx1_ASAP7_75t_R register___U2596 ( .A(register__n13349), .Y(register__n715) );
  AO22x1_ASAP7_75t_R register___U2597 ( .A1(register__net139860), .A2(register__n1603), .B1(register__n719), .B2(register__n3022), 
        .Y(register__n718) );
  CKINVDCx20_ASAP7_75t_R register___U2598 ( .A(register__n9511), .Y(register__n719) );
  INVx3_ASAP7_75t_R register___U2599 ( .A(register__net139860), .Y(register__net64688) );
  BUFx12_ASAP7_75t_R register___U2600 ( .A(register__net145247), .Y(register__net145246) );
  NOR2xp33_ASAP7_75t_R register___U2601 ( .A(register__n2002), .B(register__n6219), .Y(register__n720) );
  NOR3xp33_ASAP7_75t_R register___U2602 ( .A(register__n720), .B(register__n721), .C(register__n722), .Y(register__n10551) );
  HB1xp67_ASAP7_75t_R register___U2603 ( .A(register__n10556), .Y(register__n6219) );
  BUFx3_ASAP7_75t_R register___U2604 ( .A(register__n11182), .Y(register__n6983) );
  HB1xp67_ASAP7_75t_R register___U2605 ( .A(register__n10551), .Y(register__n5458) );
  HB1xp67_ASAP7_75t_R register___U2606 ( .A(register__n12917), .Y(register__n2951) );
  BUFx4f_ASAP7_75t_R register___U2607 ( .A(register__net103248), .Y(register__net92027) );
  BUFx4f_ASAP7_75t_R register___U2608 ( .A(register__net103248), .Y(register__net63290) );
  INVx2_ASAP7_75t_R register___U2609 ( .A(register__net63290), .Y(register__net63256) );
  HB1xp67_ASAP7_75t_R register___U2610 ( .A(register__n12759), .Y(register__n3885) );
  INVxp67_ASAP7_75t_R register___U2611 ( .A(register__n11892), .Y(register__n1635) );
  BUFx3_ASAP7_75t_R register___U2612 ( .A(RegWrite), .Y(register__n5049) );
  OAI22xp33_ASAP7_75t_R register___U2613 ( .A1(register__n12144), .A2(register__n1408), .B1(register__n8115), .B2(
        n11752), .Y(register__n723) );
  NOR2x1p5_ASAP7_75t_R register___U2614 ( .A(register__net61369), .B(register__net64052), .Y(register__n2134) );
  BUFx3_ASAP7_75t_R register___U2615 ( .A(register__n3456), .Y(register__n3043) );
  BUFx6f_ASAP7_75t_R register___U2616 ( .A(register__n11812), .Y(register__n3456) );
  NAND2xp5_ASAP7_75t_R register___U2617 ( .A(register__n1238), .B(register__n4036), .Y(register__n1088) );
  INVx1_ASAP7_75t_R register___U2618 ( .A(register__n12765), .Y(register__n725) );
  BUFx12f_ASAP7_75t_R register___U2619 ( .A(register__n1872), .Y(register__n1800) );
  HB1xp67_ASAP7_75t_R register___U2620 ( .A(register__n11779), .Y(register__n11771) );
  BUFx2_ASAP7_75t_R register___U2621 ( .A(register__n11778), .Y(register__n11769) );
  AO22x1_ASAP7_75t_R register___U2622 ( .A1(register__n9748), .A2(register__net131160), .B1(register__n10108), .B2(register__n326), .Y(register__n10773) );
  BUFx6f_ASAP7_75t_R register___U2623 ( .A(register__n2854), .Y(register__n2966) );
  INVxp67_ASAP7_75t_R register___U2624 ( .A(register__n4068), .Y(register__n6127) );
  HB1xp67_ASAP7_75t_R register___U2625 ( .A(register__n4069), .Y(register__n4068) );
  INVx6_ASAP7_75t_R register___U2626 ( .A(write_data[26]), .Y(register__n12419) );
  INVx2_ASAP7_75t_R register___U2627 ( .A(register__n1374), .Y(register__n6265) );
  NAND2xp33_ASAP7_75t_R register___U2628 ( .A(register__n727), .B(register__n1851), .Y(register__n728) );
  INVxp33_ASAP7_75t_R register___U2629 ( .A(register__net64780), .Y(register__n727) );
  INVxp67_ASAP7_75t_R register___U2630 ( .A(IF_ID_rs1[1]), .Y(register__n11132) );
  INVx6_ASAP7_75t_R register___U2631 ( .A(register__n11746), .Y(register__n1408) );
  INVx1_ASAP7_75t_R register___U2632 ( .A(register__n7577), .Y(register__n832) );
  HB1xp67_ASAP7_75t_R register___U2633 ( .A(register__n7117), .Y(register__n7116) );
  HB1xp67_ASAP7_75t_R register___U2634 ( .A(register__n4506), .Y(register__n4505) );
  INVxp33_ASAP7_75t_R register___U2635 ( .A(register__n4851), .Y(register__n808) );
  INVxp33_ASAP7_75t_R register___U2636 ( .A(register__n4851), .Y(register__n807) );
  AOI22xp5_ASAP7_75t_R register___U2637 ( .A1(register__net63212), .A2(register__n1603), .B1(register__n730), .B2(register__n3022), .Y(register__n12696) );
  CKINVDCx20_ASAP7_75t_R register___U2638 ( .A(register__net94176), .Y(register__n730) );
  HB1xp67_ASAP7_75t_R register___U2639 ( .A(register__n3743), .Y(register__n3742) );
  INVx1_ASAP7_75t_R register___U2640 ( .A(register__n1784), .Y(register__n1631) );
  INVx1_ASAP7_75t_R register___U2641 ( .A(register__n1783), .Y(register__n1784) );
  BUFx12f_ASAP7_75t_R register___U2642 ( .A(register__n3507), .Y(register__n12247) );
  BUFx6f_ASAP7_75t_R register___U2643 ( .A(register__n12247), .Y(register__n3732) );
  OAI21xp33_ASAP7_75t_R register___U2644 ( .A1(register__n2658), .A2(register__n1247), .B(register__n2681), .Y(register__n2682)
         );
  HB1xp67_ASAP7_75t_R register___U2645 ( .A(register__n11838), .Y(register__n11842) );
  HB1xp67_ASAP7_75t_R register___U2646 ( .A(register__n13237), .Y(register__n4518) );
  AND2x2_ASAP7_75t_R register___U2647 ( .A(register__C6422_net59540), .B(register__n10824), .Y(register__n798) );
  INVx3_ASAP7_75t_R register___U2648 ( .A(register__n10824), .Y(register__n8587) );
  INVx1_ASAP7_75t_R register___U2649 ( .A(register__n12588), .Y(register__n735) );
  HB1xp67_ASAP7_75t_R register___U2650 ( .A(register__n861), .Y(register__net147584) );
  HB1xp67_ASAP7_75t_R register___U2651 ( .A(register__n13317), .Y(register__n5012) );
  BUFx2_ASAP7_75t_R register___U2652 ( .A(register__n6019), .Y(register__n6018) );
  AND4x1_ASAP7_75t_R register___U2653 ( .A(register__n7607), .B(register__n124), .C(register__n7608), .D(register__n5629), .Y(
        n11078) );
  AND2x4_ASAP7_75t_R register___U2654 ( .A(rs2[4]), .B(rs2[3]), 
        .Y(register__n739) );
  INVxp67_ASAP7_75t_R register___U2655 ( .A(register__n5009), .Y(register__n6203) );
  HB1xp67_ASAP7_75t_R register___U2656 ( .A(register__n5010), .Y(register__n5009) );
  HB1xp67_ASAP7_75t_R register___U2657 ( .A(register__n2920), .Y(register__n2919) );
  HB1xp67_ASAP7_75t_R register___U2658 ( .A(register__n13223), .Y(register__n4141) );
  BUFx2_ASAP7_75t_R register___U2659 ( .A(register__n1643), .Y(register__n3832) );
  INVx1_ASAP7_75t_R register___U2660 ( .A(register__n3690), .Y(register__n1526) );
  INVx6_ASAP7_75t_R register___U2661 ( .A(register__n6465), .Y(register__n2005) );
  XNOR2xp5_ASAP7_75t_R register___U2662 ( .A(register__n11846), .B(register__n717), .Y(register__n12513) );
  INVx1_ASAP7_75t_R register___U2663 ( .A(register__net63280), .Y(register__net63248) );
  BUFx6f_ASAP7_75t_R register___U2664 ( .A(register__n12190), .Y(register__n3845) );
  HB1xp67_ASAP7_75t_R register___U2665 ( .A(register__n12996), .Y(register__n3590) );
  BUFx2_ASAP7_75t_R register___U2666 ( .A(register__n3020), .Y(register__n2969) );
  BUFx6f_ASAP7_75t_R register___U2667 ( .A(register__n2964), .Y(register__n2962) );
  INVxp67_ASAP7_75t_R register___U2668 ( .A(register__n5079), .Y(register__n6727) );
  HB1xp67_ASAP7_75t_R register___U2669 ( .A(register__n5080), .Y(register__n5079) );
  BUFx2_ASAP7_75t_R register___U2670 ( .A(register__net122408), .Y(register__net63284) );
  AND3x1_ASAP7_75t_R register___U2671 ( .A(register__n2092), .B(register__n6548), .C(register__n7150), .Y(register__n11448) );
  BUFx3_ASAP7_75t_R register___U2672 ( .A(register__net63268), .Y(register__net139893) );
  INVx2_ASAP7_75t_R register___U2673 ( .A(register__n3022), .Y(register__n1590) );
  INVx4_ASAP7_75t_R register___U2674 ( .A(register__net102359), .Y(register__net105510) );
  INVx4_ASAP7_75t_R register___U2675 ( .A(register__net137800), .Y(register__n1677) );
  HB1xp67_ASAP7_75t_R register___U2676 ( .A(register__n13219), .Y(register__n3660) );
  HB1xp67_ASAP7_75t_R register___U2677 ( .A(register__n12672), .Y(register__n7117) );
  HB1xp67_ASAP7_75t_R register___U2678 ( .A(register__n13328), .Y(register__n4069) );
  INVxp67_ASAP7_75t_R register___U2679 ( .A(register__n3220), .Y(register__n4382) );
  HB1xp67_ASAP7_75t_R register___U2680 ( .A(register__n3221), .Y(register__n3220) );
  INVx1_ASAP7_75t_R register___U2681 ( .A(register__n12895), .Y(register__n737) );
  INVx4_ASAP7_75t_R register___U2682 ( .A(register__n11816), .Y(register__n1604) );
  INVx4_ASAP7_75t_R register___U2683 ( .A(register__n2965), .Y(register__n3072) );
  INVx2_ASAP7_75t_R register___U2684 ( .A(register__n2965), .Y(register__n2950) );
  INVx1_ASAP7_75t_R register___U2685 ( .A(register__n2965), .Y(register__n1598) );
  INVx1_ASAP7_75t_R register___U2686 ( .A(register__n12929), .Y(register__n738) );
  BUFx12f_ASAP7_75t_R register___U2687 ( .A(register__n11750), .Y(register__n11746) );
  OAI22xp5_ASAP7_75t_R register___U2688 ( .A1(register__net66308), .A2(register__n7888), .B1(register__n12138), .B2(
        n1687), .Y(read_reg_data_2[12]) );
  BUFx4f_ASAP7_75t_R register___U2689 ( .A(register__net63268), .Y(register__net141048) );
  HB1xp67_ASAP7_75t_R register___U2690 ( .A(register__n12811), .Y(register__n3221) );
  INVxp67_ASAP7_75t_R register___U2691 ( .A(register__n4994), .Y(register__n6828) );
  AOI22xp5_ASAP7_75t_R register___U2692 ( .A1(register__net63284), .A2(register__n1723), .B1(register__n741), .B2(register__n1718), .Y(register__n13245) );
  CKINVDCx20_ASAP7_75t_R register___U2693 ( .A(register__net89049), .Y(register__n741) );
  CKINVDCx5p33_ASAP7_75t_R register___U2694 ( .A(register__net63284), .Y(register__net63240) );
  NOR2xp33_ASAP7_75t_R register___U2695 ( .A(register__n158), .B(register__n2387), .Y(register__n2388) );
  INVxp67_ASAP7_75t_R register___U2696 ( .A(register__n13184), .Y(register__n8240) );
  BUFx12f_ASAP7_75t_R register___U2697 ( .A(register__n11939), .Y(register__n3595) );
  BUFx6f_ASAP7_75t_R register___U2698 ( .A(register__n11948), .Y(register__n11947) );
  INVx6_ASAP7_75t_R register___U2699 ( .A(write_data[0]), .Y(register__n11948) );
  AOI22xp33_ASAP7_75t_R register___U2700 ( .A1(register__net63286), .A2(register__n473), .B1(register__n742), .B2(register__n459), 
        .Y(register__n12925) );
  CKINVDCx20_ASAP7_75t_R register___U2701 ( .A(register__net112347), .Y(register__n742) );
  AND2x2_ASAP7_75t_R register___U2702 ( .A(register__n8577), .B(register__n743), .Y(register__n10838) );
  AND2x4_ASAP7_75t_R register___U2703 ( .A(register__n11153), .B(register__n885), .Y(register__n11152) );
  AOI22xp33_ASAP7_75t_R register___U2704 ( .A1(register__n11944), .A2(register__n1584), .B1(register__n745), .B2(register__n2935), 
        .Y(register__n12717) );
  CKINVDCx20_ASAP7_75t_R register___U2705 ( .A(register__n9457), .Y(register__n745) );
  INVxp33_ASAP7_75t_R register___U2706 ( .A(register__n11944), .Y(register__n11932) );
  INVx2_ASAP7_75t_R register___U2707 ( .A(register__n3022), .Y(register__n1584) );
  CKINVDCx20_ASAP7_75t_R register___U2708 ( .A(register__n12516), .Y(register__n746) );
  INVx1_ASAP7_75t_R register___U2709 ( .A(register__n12521), .Y(register__n6759) );
  AND2x4_ASAP7_75t_R register___U2710 ( .A(register__n149), .B(register__n7020), .Y(register__C6423_net60466) );
  HB1xp67_ASAP7_75t_R register___U2711 ( .A(register__n13315), .Y(register__n4506) );
  INVx1_ASAP7_75t_R register___U2712 ( .A(register__n2936), .Y(register__n1596) );
  INVx1_ASAP7_75t_R register___U2713 ( .A(register__n12075), .Y(register__n12062) );
  AND2x4_ASAP7_75t_R register___U2714 ( .A(register__n1476), .B(register__n1513), .Y(register__n8752) );
  INVx2_ASAP7_75t_R register___U2715 ( .A(register__n3184), .Y(register__n1309) );
  HB1xp67_ASAP7_75t_R register___U2716 ( .A(register__n13213), .Y(register__n4143) );
  INVx3_ASAP7_75t_R register___U2717 ( .A(register__n4641), .Y(register__n11754) );
  INVx1_ASAP7_75t_R register___U2718 ( .A(register__n12493), .Y(register__n748) );
  AND2x2_ASAP7_75t_R register___U2719 ( .A(register__n12492), .B(register__n830), .Y(register__n12493) );
  OAI22xp5_ASAP7_75t_R register___U2720 ( .A1(register__n54), .A2(register__n7324), .B1(register__net61369), .B2(register__n12206), .Y(read_reg_data_1[16]) );
  AND2x2_ASAP7_75t_R register___U2721 ( .A(register__n11720), .B(register__n1953), .Y(register__n1966) );
  INVx2_ASAP7_75t_R register___U2722 ( .A(register__n3072), .Y(register__n11894) );
  OAI22xp33_ASAP7_75t_R register___U2723 ( .A1(register__n12251), .A2(register__n1408), .B1(register__net89877), .B2(
        n2886), .Y(register__n749) );
  INVxp67_ASAP7_75t_R register___U2724 ( .A(register__n3926), .Y(register__n7078) );
  HB1xp67_ASAP7_75t_R register___U2725 ( .A(register__n3927), .Y(register__n3926) );
  NOR2xp67_ASAP7_75t_R register___U2726 ( .A(register__n10210), .B(register__n11799), .Y(register__n1170) );
  BUFx12f_ASAP7_75t_R register___U2727 ( .A(register__n3564), .Y(register__n11799) );
  INVx3_ASAP7_75t_R register___U2728 ( .A(register__net63286), .Y(register__net63252) );
  INVxp33_ASAP7_75t_R register___U2729 ( .A(register__n1137), .Y(register__n1151) );
  INVx1_ASAP7_75t_R register___U2730 ( .A(register__n103), .Y(register__n1146) );
  INVxp67_ASAP7_75t_R register___U2731 ( .A(register__n103), .Y(register__n1148) );
  INVxp67_ASAP7_75t_R register___U2732 ( .A(register__n103), .Y(register__n1150) );
  INVx1_ASAP7_75t_R register___U2733 ( .A(register__n103), .Y(register__n1147) );
  INVxp33_ASAP7_75t_R register___U2734 ( .A(register__n103), .Y(register__n1149) );
  OR2x2_ASAP7_75t_R register___U2735 ( .A(register__n48), .B(register__n9178), .Y(register__n751) );
  OR2x2_ASAP7_75t_R register___U2736 ( .A(register__net61369), .B(register__net63216), .Y(register__n752) );
  AO211x2_ASAP7_75t_R register___U2737 ( .A1(register__net89689), .A2(register__n366), .B(register__n753), .C(register__n754), 
        .Y(register__n2411) );
  AO21x1_ASAP7_75t_R register___U2738 ( .A1(register__net120788), .A2(register__net90965), .B(register__n2393), .Y(register__n753) );
  INVxp33_ASAP7_75t_R register___U2739 ( .A(register__n7087), .Y(register__n1525) );
  INVx1_ASAP7_75t_R register___U2740 ( .A(register__n12583), .Y(register__n755) );
  AO22x1_ASAP7_75t_R register___U2741 ( .A1(register__net90905), .A2(register__net109849), .B1(register__net89997), 
        .B2(register__C6423_net61348), .Y(register__n11296) );
  HB1xp67_ASAP7_75t_R register___U2742 ( .A(register__n11385), .Y(register__n3246) );
  AO22x1_ASAP7_75t_R register___U2743 ( .A1(register__n9658), .A2(register__net109849), .B1(register__n9985), .B2(
        C6423_net61348), .Y(register__n11173) );
  INVx2_ASAP7_75t_R register___U2744 ( .A(register__n1136), .Y(register__n1143) );
  AO22x1_ASAP7_75t_R register___U2745 ( .A1(register__n10497), .A2(register__net129747), .B1(register__n8787), .B2(
        C6422_net70296), .Y(register__n10562) );
  AO22x1_ASAP7_75t_R register___U2746 ( .A1(register__net103466), .A2(register__C6422_net60422), .B1(register__net89461), .B2(register__net123857), .Y(register__n10709) );
  AO22x1_ASAP7_75t_R register___U2747 ( .A1(register__n9762), .A2(register__C6422_net60422), .B1(register__n10155), 
        .B2(register__net123857), .Y(register__n10648) );
  BUFx3_ASAP7_75t_R register___U2748 ( .A(register__n5410), .Y(register__n5409) );
  BUFx2_ASAP7_75t_R register___U2749 ( .A(register__n5415), .Y(register__n5414) );
  INVx1_ASAP7_75t_R register___U2750 ( .A(register__n12570), .Y(register__n757) );
  INVxp67_ASAP7_75t_R register___U2751 ( .A(register__n4445), .Y(register__n6702) );
  AO22x1_ASAP7_75t_R register___U2752 ( .A1(register__n9266), .A2(register__net117658), .B1(register__n10319), .B2(register__n836), .Y(register__n10848) );
  AO22x1_ASAP7_75t_R register___U2753 ( .A1(register__n9573), .A2(register__net117658), .B1(register__n9429), .B2(register__n834), 
        .Y(register__n10827) );
  AO22x1_ASAP7_75t_R register___U2754 ( .A1(register__n9252), .A2(register__net117658), .B1(register__n10056), .B2(register__n834), .Y(register__n10917) );
  AO22x1_ASAP7_75t_R register___U2755 ( .A1(register__net93805), .A2(register__C6422_net60408), .B1(register__net103457), .B2(register__n836), .Y(register__n10704) );
  AO22x1_ASAP7_75t_R register___U2756 ( .A1(register__n9248), .A2(register__net117658), .B1(register__n10052), .B2(register__n842), .Y(register__n10961) );
  AO22x1_ASAP7_75t_R register___U2757 ( .A1(register__n9250), .A2(register__net117658), .B1(register__n7458), .B2(register__n834), 
        .Y(register__n10938) );
  NOR2xp33_ASAP7_75t_R register___U2758 ( .A(register__n1995), .B(register__n5728), .Y(register__n759) );
  NOR2xp33_ASAP7_75t_R register___U2759 ( .A(register__n1800), .B(register__n6214), .Y(register__n760) );
  HB1xp67_ASAP7_75t_R register___U2760 ( .A(register__n11503), .Y(register__n5728) );
  HB1xp67_ASAP7_75t_R register___U2761 ( .A(register__n11504), .Y(register__n6214) );
  AND2x2_ASAP7_75t_R register___U2762 ( .A(register__n12495), .B(register__n796), .Y(register__n12500) );
  INVx6_ASAP7_75t_R register___U2763 ( .A(register__n108), .Y(register__n12171) );
  HB1xp67_ASAP7_75t_R register___U2764 ( .A(register__n667), .Y(register__net63268) );
  HB1xp67_ASAP7_75t_R register___U2765 ( .A(register__net63268), .Y(register__net63276) );
  INVx2_ASAP7_75t_R register___U2766 ( .A(register__net63282), .Y(register__net63250) );
  INVx2_ASAP7_75t_R register___U2767 ( .A(register__net73055), .Y(register__n2105) );
  BUFx12_ASAP7_75t_R register___U2768 ( .A(register__n3646), .Y(register__n3838) );
  HB1xp67_ASAP7_75t_R register___U2769 ( .A(register__n13110), .Y(register__n3927) );
  AOI21xp5_ASAP7_75t_R register___U2770 ( .A1(register__net134749), .A2(register__net93717), .B(register__n2680), .Y(
        n2681) );
  NOR3x1_ASAP7_75t_R register___U2771 ( .A(register__n7958), .B(register__n7957), .C(register__n7956), .Y(register__n763) );
  BUFx6f_ASAP7_75t_R register___U2772 ( .A(register__n3071), .Y(register__n2970) );
  INVxp67_ASAP7_75t_R register___U2773 ( .A(register__n2118), .Y(register__n2121) );
  AO22x1_ASAP7_75t_R register___U2774 ( .A1(register__n9887), .A2(register__n3), .B1(register__n10311), .B2(register__n233), .Y(
        n10858) );
  HB1xp67_ASAP7_75t_R register___U2775 ( .A(register__n4995), .Y(register__n4994) );
  AO22x1_ASAP7_75t_R register___U2776 ( .A1(register__net90229), .A2(register__n413), .B1(register__net89005), .B2(
        net126602), .Y(register__n11086) );
  AO22x1_ASAP7_75t_R register___U2777 ( .A1(register__n9640), .A2(register__n413), .B1(register__n9951), .B2(
        C6422_net60401), .Y(register__n10536) );
  AO22x1_ASAP7_75t_R register___U2778 ( .A1(register__n10432), .A2(register__n413), .B1(register__n10428), .B2(
        net126602), .Y(register__n10686) );
  AO22x1_ASAP7_75t_R register___U2779 ( .A1(register__n8759), .A2(register__n413), .B1(register__n9945), .B2(register__net126602), 
        .Y(register__n10939) );
  AND2x4_ASAP7_75t_R register___U2780 ( .A(register__n11719), .B(register__n389), .Y(register__C6423_net61325) );
  BUFx4f_ASAP7_75t_R register___U2781 ( .A(register__n4122), .Y(register__n2936) );
  BUFx3_ASAP7_75t_R register___U2782 ( .A(register__n11796), .Y(register__n11791) );
  AO22x1_ASAP7_75t_R register___U2783 ( .A1(register__n6286), .A2(register__n413), .B1(register__n4757), .B2(register__net126602), 
        .Y(register__n10962) );
  INVx1_ASAP7_75t_R register___U2784 ( .A(register__n10862), .Y(register__n764) );
  INVx6_ASAP7_75t_R register___U2785 ( .A(register__n3190), .Y(register__n3071) );
  NAND3xp33_ASAP7_75t_R register___U2786 ( .A(register__n10717), .B(register__n10716), .C(register__n1021), .Y(register__n2216)
         );
  NOR2xp33_ASAP7_75t_R register___U2787 ( .A(register__n765), .B(register__n766), .Y(register__n11522) );
  BUFx3_ASAP7_75t_R register___U2788 ( .A(register__n11526), .Y(register__n7867) );
  HB1xp67_ASAP7_75t_R register___U2789 ( .A(register__n11522), .Y(register__n5804) );
  AND2x2_ASAP7_75t_R register___U2790 ( .A(register__n5441), .B(register__n7052), .Y(register__n7996) );
  AOI21xp33_ASAP7_75t_R register___U2791 ( .A1(register__n326), .A2(register__net89645), .B(register__n2674), .Y(register__n2675)
         );
  INVx4_ASAP7_75t_R register___U2792 ( .A(register__n11554), .Y(register__n1570) );
  BUFx6f_ASAP7_75t_R register___U2793 ( .A(register__net64900), .Y(register__net64896) );
  BUFx6f_ASAP7_75t_R register___U2794 ( .A(register__C6423_net61331), .Y(register__n2025) );
  INVx4_ASAP7_75t_R register___U2795 ( .A(register__n2023), .Y(register__n2024) );
  BUFx6f_ASAP7_75t_R register___U2796 ( .A(register__n2024), .Y(register__net130032) );
  INVx6_ASAP7_75t_R register___U2797 ( .A(register__n2025), .Y(register__n2023) );
  INVx6_ASAP7_75t_R register___U2798 ( .A(register__net130032), .Y(register__net130031) );
  BUFx6f_ASAP7_75t_R register___U2799 ( .A(register__net130031), .Y(register__net99861) );
  HB1xp67_ASAP7_75t_R register___U2800 ( .A(register__net99861), .Y(register__net130030) );
  INVx1_ASAP7_75t_R register___U2801 ( .A(register__n1136), .Y(register__n1142) );
  INVx2_ASAP7_75t_R register___U2802 ( .A(register__n1136), .Y(register__n1145) );
  HB1xp67_ASAP7_75t_R register___U2803 ( .A(register__n13226), .Y(register__n5579) );
  INVx1_ASAP7_75t_R register___U2804 ( .A(register__n13268), .Y(register__n3871) );
  INVx2_ASAP7_75t_R register___U2805 ( .A(register__n11367), .Y(register__n1047) );
  CKINVDCx8_ASAP7_75t_R register___U2806 ( .A(register__net137417), .Y(register__net122250) );
  NOR3xp33_ASAP7_75t_R register___U2807 ( .A(register__n2604), .B(register__n2625), .C(register__n2626), .Y(register__n2624) );
  OAI22xp5_ASAP7_75t_R register___U2808 ( .A1(register__net66320), .A2(register__n7941), .B1(register__net62710), .B2(
        n1687), .Y(read_reg_data_2[31]) );
  INVxp67_ASAP7_75t_R register___U2809 ( .A(register__n11894), .Y(register__n1602) );
  INVx6_ASAP7_75t_R register___U2810 ( .A(register__n3439), .Y(register__n12054) );
  INVx2_ASAP7_75t_R register___U2811 ( .A(register__net127289), .Y(register__n1684) );
  INVx3_ASAP7_75t_R register___U2812 ( .A(IF_ID_rs1[2]), .Y(register__n1513) );
  BUFx6f_ASAP7_75t_R register___U2813 ( .A(register__n4850), .Y(register__n3190) );
  BUFx6f_ASAP7_75t_R register___U2814 ( .A(register__C6423_net68516), .Y(register__net107120) );
  INVxp67_ASAP7_75t_R register___U2815 ( .A(register__n5331), .Y(register__n9220) );
  HB1xp67_ASAP7_75t_R register___U2816 ( .A(register__n12647), .Y(register__n4396) );
  NOR3x1_ASAP7_75t_R register___U2817 ( .A(register__n74), .B(register__n226), .C(register__n4921), .Y(register__n7324) );
  HB1xp67_ASAP7_75t_R register___U2818 ( .A(register__n6419), .Y(register__n4558) );
  INVxp33_ASAP7_75t_R register___U2819 ( .A(register__n4556), .Y(register__n6419) );
  AOI22xp33_ASAP7_75t_R register___U2820 ( .A1(register__net145264), .A2(register__n1972), .B1(register__n1130), .B2(
        n1131), .Y(register__n12914) );
  AOI21xp5_ASAP7_75t_R register___U2821 ( .A1(register__n39), .A2(register__net104596), .B(register__n2352), .Y(register__n2354)
         );
  NOR2xp67_ASAP7_75t_R register___U2822 ( .A(register__n2356), .B(register__n2335), .Y(register__n2355) );
  HB1xp67_ASAP7_75t_R register___U2823 ( .A(register__n10587), .Y(register__n4445) );
  BUFx6f_ASAP7_75t_R register___U2824 ( .A(register__net144708), .Y(register__net64816) );
  INVx1_ASAP7_75t_R register___U2825 ( .A(register__n2011), .Y(register__n1918) );
  INVx4_ASAP7_75t_R register___U2826 ( .A(register__n11877), .Y(register__n2010) );
  INVx4_ASAP7_75t_R register___U2827 ( .A(register__n3309), .Y(register__n2285) );
  NOR4xp75_ASAP7_75t_R register___U2828 ( .A(register__n1896), .B(register__n2544), .C(register__n2539), .D(register__n2542), .Y(
        n2568) );
  NOR2x1p5_ASAP7_75t_R register___U2829 ( .A(register__n112), .B(register__n2543), .Y(register__n2544) );
  INVxp67_ASAP7_75t_R register___U2830 ( .A(register__n2019), .Y(register__n769) );
  INVx1_ASAP7_75t_R register___U2831 ( .A(register__n2019), .Y(register__n770) );
  INVxp67_ASAP7_75t_R register___U2832 ( .A(register__net150876), .Y(register__net150890) );
  INVxp67_ASAP7_75t_R register___U2833 ( .A(register__net150880), .Y(register__net150892) );
  INVx5_ASAP7_75t_R register___U2834 ( .A(register__n2019), .Y(register__net150889) );
  INVx4_ASAP7_75t_R register___U2835 ( .A(register__n1905), .Y(register__n1906) );
  INVx2_ASAP7_75t_R register___U2836 ( .A(register__net150889), .Y(register__n1905) );
  INVx1_ASAP7_75t_R register___U2837 ( .A(register__n10735), .Y(register__n771) );
  INVxp67_ASAP7_75t_R register___U2838 ( .A(write_data[25]), .Y(register__net63222) );
  INVxp67_ASAP7_75t_R register___U2839 ( .A(register__n13139), .Y(register__n4049) );
  BUFx6f_ASAP7_75t_R register___U2840 ( .A(register__n8564), .Y(register__n8562) );
  INVx2_ASAP7_75t_R register___U2841 ( .A(register__n4932), .Y(register__n7958) );
  OA22x2_ASAP7_75t_R register___U2842 ( .A1(register__n12083), .A2(register__n11868), .B1(register__n6626), .B2(register__n2886), 
        .Y(register__n13278) );
  BUFx4_ASAP7_75t_R register___U2843 ( .A(register__n8356), .Y(register__n6626) );
  BUFx12f_ASAP7_75t_R register___U2844 ( .A(register__n4475), .Y(register__n11739) );
  CKINVDCx5p33_ASAP7_75t_R register___U2845 ( .A(register__net62700), .Y(register__net62666) );
  INVxp67_ASAP7_75t_R register___U2846 ( .A(register__n1937), .Y(register__n1934) );
  INVxp67_ASAP7_75t_R register___U2847 ( .A(register__n2814), .Y(register__n1941) );
  INVx1_ASAP7_75t_R register___U2848 ( .A(register__n2005), .Y(register__n2007) );
  INVx1_ASAP7_75t_R register___U2849 ( .A(register__n2005), .Y(register__n2009) );
  INVx1_ASAP7_75t_R register___U2850 ( .A(register__n2005), .Y(register__n2006) );
  AO22x1_ASAP7_75t_R register___U2851 ( .A1(register__net90521), .A2(register__n3), .B1(register__net89397), .B2(register__n281), 
        .Y(register__n10817) );
  AO22x1_ASAP7_75t_R register___U2852 ( .A1(register__n10442), .A2(register__n1909), .B1(register__n10426), .B2(register__n381), 
        .Y(register__n11054) );
  AO22x1_ASAP7_75t_R register___U2853 ( .A1(register__n9652), .A2(register__n1909), .B1(register__n9979), .B2(register__n381), 
        .Y(register__n10610) );
  INVx1_ASAP7_75t_R register___U2854 ( .A(register__n1363), .Y(register__n13307) );
  INVx1_ASAP7_75t_R register___U2855 ( .A(register__n13199), .Y(register__n776) );
  INVx4_ASAP7_75t_R register___U2856 ( .A(register__n3338), .Y(register__n11868) );
  BUFx3_ASAP7_75t_R register___U2857 ( .A(register__n10658), .Y(register__n4933) );
  HB1xp67_ASAP7_75t_R register___U2858 ( .A(register__n4924), .Y(register__n4923) );
  BUFx12f_ASAP7_75t_R register___U2859 ( .A(register__n12384), .Y(register__n12388) );
  HB1xp67_ASAP7_75t_R register___U2860 ( .A(register__n3282), .Y(register__n3263) );
  BUFx3_ASAP7_75t_R register___U2861 ( .A(register__net122250), .Y(register__net122247) );
  INVx1_ASAP7_75t_R register___U2862 ( .A(register__n12709), .Y(register__n777) );
  AND2x2_ASAP7_75t_R register___U2863 ( .A(register__n778), .B(register__n8314), .Y(register__n8645) );
  INVx4_ASAP7_75t_R register___U2864 ( .A(register__net64458), .Y(register__net64426) );
  INVx1_ASAP7_75t_R register___U2865 ( .A(register__n11013), .Y(register__n779) );
  HB1xp67_ASAP7_75t_R register___U2866 ( .A(register__n12634), .Y(register__n4510) );
  HB1xp67_ASAP7_75t_R register___U2867 ( .A(register__n12613), .Y(register__n4534) );
  OA22x2_ASAP7_75t_R register___U2868 ( .A1(register__n781), .A2(register__n11868), .B1(register__n10307), .B2(register__n3338), 
        .Y(register__n780) );
  INVxp67_ASAP7_75t_R register___U2869 ( .A(register__n11271), .Y(register__n782) );
  BUFx6f_ASAP7_75t_R register___U2870 ( .A(register__n3535), .Y(register__n3594) );
  OAI211xp5_ASAP7_75t_R register___U2871 ( .A1(register__n1507), .A2(register__n2246), .B(register__n12508), .C(register__n2053), 
        .Y(register__n783) );
  AO22x1_ASAP7_75t_R register___U2872 ( .A1(register__n9654), .A2(register__n156), .B1(register__n9981), .B2(register__n233), .Y(
        n10587) );
  INVx1_ASAP7_75t_R register___U2873 ( .A(register__n11552), .Y(register__n784) );
  NOR2xp33_ASAP7_75t_R register___U2874 ( .A(register__n2081), .B(register__n6763), .Y(register__n785) );
  HB1xp67_ASAP7_75t_R register___U2875 ( .A(register__n11063), .Y(register__n6763) );
  HB1xp67_ASAP7_75t_R register___U2876 ( .A(register__n11065), .Y(register__n6473) );
  INVx1_ASAP7_75t_R register___U2877 ( .A(register__n12690), .Y(register__n788) );
  INVx2_ASAP7_75t_R register___U2878 ( .A(register__n8274), .Y(register__n1479) );
  AO22x1_ASAP7_75t_R register___U2879 ( .A1(register__net63220), .A2(register__n1058), .B1(register__n790), .B2(register__n1137), 
        .Y(register__n789) );
  CKINVDCx20_ASAP7_75t_R register___U2880 ( .A(register__net94168), .Y(register__n790) );
  HB1xp67_ASAP7_75t_R register___U2881 ( .A(register__n3342), .Y(register__n12390) );
  HB1xp67_ASAP7_75t_R register___U2882 ( .A(register__n3300), .Y(register__n12387) );
  BUFx6f_ASAP7_75t_R register___U2883 ( .A(register__n3071), .Y(register__n4122) );
  CKINVDCx10_ASAP7_75t_R register___U2884 ( .A(register__net91939), .Y(register__net64418) );
  AND2x6_ASAP7_75t_R register___U2885 ( .A(register__n12495), .B(register__n3407), .Y(register__n5720) );
  HB1xp67_ASAP7_75t_R register___U2886 ( .A(register__n3604), .Y(register__n3471) );
  BUFx6f_ASAP7_75t_R register___U2887 ( .A(register__n3471), .Y(register__n4639) );
  NOR2xp33_ASAP7_75t_R register___U2888 ( .A(register__n157), .B(register__n2655), .Y(register__n2657) );
  NOR2xp33_ASAP7_75t_R register___U2889 ( .A(register__n158), .B(register__n2339), .Y(register__n2340) );
  AO22x1_ASAP7_75t_R register___U2890 ( .A1(register__n9333), .A2(register__n3), .B1(register__n8789), .B2(register__n281), .Y(
        n10837) );
  AOI22xp33_ASAP7_75t_R register___U2891 ( .A1(register__net64458), .A2(register__n5721), .B1(register__n791), .B2(
        n1411), .Y(register__n12999) );
  CKINVDCx20_ASAP7_75t_R register___U2892 ( .A(register__net90393), .Y(register__n791) );
  CKINVDCx5p33_ASAP7_75t_R register___U2893 ( .A(register__n1411), .Y(register__n1418) );
  HB1xp67_ASAP7_75t_R register___U2894 ( .A(register__n5442), .Y(register__n12218) );
  HB1xp67_ASAP7_75t_R register___U2895 ( .A(register__n3667), .Y(register__n12220) );
  BUFx2_ASAP7_75t_R register___U2896 ( .A(register__net143491), .Y(register__net63034) );
  HB1xp67_ASAP7_75t_R register___U2897 ( .A(register__n3359), .Y(register__n4843) );
  BUFx6f_ASAP7_75t_R register___U2898 ( .A(register__n5353), .Y(register__n3475) );
  INVxp33_ASAP7_75t_R register___U2899 ( .A(register__net106927), .Y(register__n1204) );
  INVxp33_ASAP7_75t_R register___U2900 ( .A(register__net106927), .Y(register__n2151) );
  OAI22xp33_ASAP7_75t_R register___U2901 ( .A1(register__net64922), .A2(register__n11861), .B1(register__n10044), .B2(
        n1161), .Y(register__n792) );
  INVxp33_ASAP7_75t_R register___U2902 ( .A(register__net122579), .Y(register__n793) );
  INVxp67_ASAP7_75t_R register___U2903 ( .A(register__n11444), .Y(register__n794) );
  BUFx12f_ASAP7_75t_R register___U2904 ( .A(register__n12222), .Y(register__n3645) );
  INVx1_ASAP7_75t_R register___U2905 ( .A(register__n12625), .Y(register__n795) );
  BUFx6f_ASAP7_75t_R register___U2906 ( .A(register__net136186), .Y(register__net63052) );
  AO22x1_ASAP7_75t_R register___U2907 ( .A1(register__net91033), .A2(register__n128), .B1(register__net89865), .B2(
        n1443), .Y(register__n11287) );
  BUFx12f_ASAP7_75t_R register___U2908 ( .A(register__n3571), .Y(register__n3727) );
  BUFx2_ASAP7_75t_R register___U2909 ( .A(register__n12336), .Y(register__n8244) );
  BUFx6f_ASAP7_75t_R register___U2910 ( .A(register__n8244), .Y(register__n3517) );
  AO22x1_ASAP7_75t_R register___U2911 ( .A1(register__n9907), .A2(register__n3), .B1(register__n10210), .B2(register__n1578), .Y(
        n10800) );
  AO22x1_ASAP7_75t_R register___U2912 ( .A1(register__n9728), .A2(register__n1909), .B1(register__n10183), .B2(register__n1578), 
        .Y(register__n10654) );
  AND4x1_ASAP7_75t_R register___U2913 ( .A(register__n8233), .B(register__n8232), .C(register__n8231), .D(register__n2900), .Y(
        n11219) );
  NOR2xp67_ASAP7_75t_R register___U2914 ( .A(register__n797), .B(register__n798), .Y(register__n10822) );
  BUFx3_ASAP7_75t_R register___U2915 ( .A(register__n10823), .Y(register__n8836) );
  HB1xp67_ASAP7_75t_R register___U2916 ( .A(register__n10822), .Y(register__n4924) );
  HB1xp67_ASAP7_75t_R register___U2917 ( .A(register__n4557), .Y(register__n4556) );
  INVx1_ASAP7_75t_R register___U2918 ( .A(register__n13308), .Y(register__n803) );
  BUFx12f_ASAP7_75t_R register___U2919 ( .A(register__net141957), .Y(register__net141956) );
  BUFx12f_ASAP7_75t_R register___U2920 ( .A(register__n3601), .Y(register__n4837) );
  HB1xp67_ASAP7_75t_R register___U2921 ( .A(register__n12393), .Y(register__n3300) );
  INVx1_ASAP7_75t_R register___U2922 ( .A(register__n13154), .Y(register__n8664) );
  INVx3_ASAP7_75t_R register___U2923 ( .A(register__n1136), .Y(register__n1144) );
  INVx2_ASAP7_75t_R register___U2924 ( .A(register__n3032), .Y(register__n1166) );
  INVx2_ASAP7_75t_R register___U2925 ( .A(register__n5319), .Y(register__n8285) );
  INVxp33_ASAP7_75t_R register___U2926 ( .A(register__n118), .Y(register__n804) );
  INVx1_ASAP7_75t_R register___U2927 ( .A(register__n12641), .Y(register__n805) );
  INVxp33_ASAP7_75t_R register___U2928 ( .A(register__n4851), .Y(register__n809) );
  INVxp33_ASAP7_75t_R register___U2929 ( .A(register__n4851), .Y(register__n810) );
  INVxp33_ASAP7_75t_R register___U2930 ( .A(register__n4851), .Y(register__n811) );
  INVxp33_ASAP7_75t_R register___U2931 ( .A(register__n4851), .Y(register__n812) );
  CKINVDCx6p67_ASAP7_75t_R register___U2932 ( .A(register__n2163), .Y(register__n1901) );
  INVx2_ASAP7_75t_R register___U2933 ( .A(register__n3867), .Y(register__n11857) );
  INVx2_ASAP7_75t_R register___U2934 ( .A(register__n3866), .Y(register__n11856) );
  AND4x1_ASAP7_75t_R register___U2935 ( .A(register__n1685), .B(register__n782), .C(register__n6056), .D(register__n4681), .Y(
        n11261) );
  HB1xp67_ASAP7_75t_R register___U2936 ( .A(register__n12717), .Y(register__n4652) );
  INVx1_ASAP7_75t_R register___U2937 ( .A(register__net74027), .Y(register__n2145) );
  INVxp33_ASAP7_75t_R register___U2938 ( .A(register__net74027), .Y(register__n1203) );
  INVx1_ASAP7_75t_R register___U2939 ( .A(register__n13269), .Y(register__n819) );
  INVxp67_ASAP7_75t_R register___U2940 ( .A(register__n733), .Y(register__n12235) );
  INVx1_ASAP7_75t_R register___U2941 ( .A(register__n12245), .Y(register__n12232) );
  AND2x2_ASAP7_75t_R register___U2942 ( .A(rs2[4]), .B(register__n1432), .Y(register__n820) );
  INVx1_ASAP7_75t_R register___U2943 ( .A(register__n13284), .Y(register__n822) );
  BUFx12f_ASAP7_75t_R register___U2944 ( .A(register__n3646), .Y(register__n12108) );
  HB1xp67_ASAP7_75t_R register___U2945 ( .A(register__n3341), .Y(register__n12385) );
  INVxp67_ASAP7_75t_R register___U2946 ( .A(register__n12970), .Y(register__n4986) );
  BUFx6f_ASAP7_75t_R register___U2947 ( .A(register__n3648), .Y(register__n3647) );
  BUFx4f_ASAP7_75t_R register___U2948 ( .A(register__n4577), .Y(register__n12274) );
  BUFx6f_ASAP7_75t_R register___U2949 ( .A(register__n4576), .Y(register__n12268) );
  BUFx3_ASAP7_75t_R register___U2950 ( .A(register__n12393), .Y(register__n12392) );
  INVx1_ASAP7_75t_R register___U2951 ( .A(register__n13283), .Y(register__n823) );
  INVx1_ASAP7_75t_R register___U2952 ( .A(register__n13274), .Y(register__n824) );
  OAI21xp33_ASAP7_75t_R register___U2953 ( .A1(register__n2552), .A2(register__n912), .B(register__n2572), .Y(register__n2571) );
  CKINVDCx10_ASAP7_75t_R register___U2954 ( .A(register__n3234), .Y(register__n7259) );
  BUFx5_ASAP7_75t_R register___U2955 ( .A(register__n3235), .Y(register__n3234) );
  INVx3_ASAP7_75t_R register___U2956 ( .A(register__n11744), .Y(register__n1409) );
  BUFx2_ASAP7_75t_R register___U2957 ( .A(register__net63276), .Y(register__net63282) );
  AND2x2_ASAP7_75t_R register___U2958 ( .A(register__n9389), .B(register__n1128), .Y(register__n830) );
  INVx3_ASAP7_75t_R register___U2959 ( .A(register__net74029), .Y(register__net123512) );
  INVx3_ASAP7_75t_R register___U2960 ( .A(register__net123512), .Y(register__net106927) );
  INVx1_ASAP7_75t_R register___U2961 ( .A(register__n13282), .Y(register__n826) );
  INVxp33_ASAP7_75t_R register___U2962 ( .A(register__net122579), .Y(register__n915) );
  AND3x1_ASAP7_75t_R register___U2963 ( .A(register__n827), .B(register__n11055), .C(register__n358), .Y(register__n9177) );
  INVx3_ASAP7_75t_R register___U2964 ( .A(register__n12269), .Y(register__n12256) );
  NOR2xp33_ASAP7_75t_R register___U2965 ( .A(register__n1800), .B(register__n6468), .Y(register__n2754) );
  OAI22xp5_ASAP7_75t_R register___U2966 ( .A1(register__n53), .A2(register__n7940), .B1(register__net61369), .B2(register__n12294), .Y(read_reg_data_1[19]) );
  INVx3_ASAP7_75t_R register___U2967 ( .A(register__n11973), .Y(register__n11957) );
  BUFx6f_ASAP7_75t_R register___U2968 ( .A(register__n7611), .Y(register__n11973) );
  HB1xp67_ASAP7_75t_R register___U2969 ( .A(register__n13316), .Y(register__n5010) );
  OAI22xp5_ASAP7_75t_R register___U2970 ( .A1(register__net66306), .A2(register__n9175), .B1(register__n12094), .B2(
        n1687), .Y(read_reg_data_2[9]) );
  INVxp67_ASAP7_75t_R register___U2971 ( .A(register__n5270), .Y(register__n8609) );
  HB1xp67_ASAP7_75t_R register___U2972 ( .A(register__n5271), .Y(register__n5270) );
  HB1xp67_ASAP7_75t_R register___U2973 ( .A(register__n5332), .Y(register__n5331) );
  BUFx6f_ASAP7_75t_R register___U2974 ( .A(register__net63286), .Y(register__net63280) );
  INVx4_ASAP7_75t_R register___U2975 ( .A(register__n3669), .Y(register__n11924) );
  INVxp67_ASAP7_75t_R register___U2976 ( .A(register__n12813), .Y(register__n4275) );
  AND2x4_ASAP7_75t_R register___U2977 ( .A(register__n12492), .B(register__n3500), .Y(register__n10517) );
  INVx1_ASAP7_75t_R register___U2978 ( .A(register__n7486), .Y(register__n1314) );
  HB1xp67_ASAP7_75t_R register___U2979 ( .A(register__n12652), .Y(register__n4406) );
  OAI21xp33_ASAP7_75t_R register___U2980 ( .A1(register__C6423_net60777), .A2(register__n1987), .B(register__n2616), 
        .Y(register__n2615) );
  INVxp67_ASAP7_75t_R register___U2981 ( .A(register__n3550), .Y(register__n5237) );
  INVx1_ASAP7_75t_R register___U2982 ( .A(register__n12659), .Y(register__n828) );
  INVx1_ASAP7_75t_R register___U2983 ( .A(register__n13112), .Y(register__n829) );
  OR2x6_ASAP7_75t_R register___U2984 ( .A(register__n6759), .B(register__n6431), .Y(register__net61369) );
  OAI22xp5_ASAP7_75t_R register___U2985 ( .A1(register__n54), .A2(register__n9177), .B1(register__net61369), .B2(register__n12436), .Y(read_reg_data_1[28]) );
  AOI222xp33_ASAP7_75t_R register___U2986 ( .A1(register__C6423_net60464), .A2(register__n10407), .B1(
        C6423_net60466), .B2(register__n9547), .C1(register__n831), .C2(register__n832), .Y(register__n11619) );
  INVx2_ASAP7_75t_R register___U2987 ( .A(write_data[22]), .Y(register__n12393) );
  BUFx6f_ASAP7_75t_R register___U2988 ( .A(register__net147583), .Y(register__net139016) );
  BUFx6f_ASAP7_75t_R register___U2989 ( .A(register__net148003), .Y(register__net100539) );
  INVx6_ASAP7_75t_R register___U2990 ( .A(register__net148409), .Y(register__net64016) );
  INVx3_ASAP7_75t_R register___U2991 ( .A(register__net63196), .Y(register__net63164) );
  INVxp67_ASAP7_75t_R register___U2992 ( .A(register__n4206), .Y(register__n6433) );
  HB1xp67_ASAP7_75t_R register___U2993 ( .A(register__n4061), .Y(register__n4060) );
  INVx1_ASAP7_75t_R register___U2994 ( .A(register__n838), .Y(register__n833) );
  INVxp67_ASAP7_75t_R register___U2995 ( .A(register__n_cell_124812_net160762), .Y(register__n840) );
  INVxp33_ASAP7_75t_R register___U2996 ( .A(register__n260), .Y(register__n842) );
  NOR2xp67_ASAP7_75t_R register___U2997 ( .A(register__n1687), .B(register__net130838), .Y(register__n2718) );
  BUFx6f_ASAP7_75t_R register___U2998 ( .A(register__net145202), .Y(register__net63196) );
  AND2x2_ASAP7_75t_R register___U2999 ( .A(register__n12183), .B(register__n9379), .Y(register__n2770) );
  BUFx3_ASAP7_75t_R register___U3000 ( .A(register__n3668), .Y(register__n3504) );
  BUFx3_ASAP7_75t_R register___U3001 ( .A(register__n3152), .Y(register__n11822) );
  AND2x2_ASAP7_75t_R register___U3002 ( .A(register__n11540), .B(register__n11541), .Y(register__n843) );
  NOR4xp25_ASAP7_75t_R register___U3003 ( .A(register__n4220), .B(register__n1228), .C(register__n11555), .D(register__n11556), 
        .Y(register__n11541) );
  BUFx12_ASAP7_75t_R register___U3004 ( .A(register__n3993), .Y(register__n12041) );
  INVxp33_ASAP7_75t_R register___U3005 ( .A(register__n3993), .Y(register__n1019) );
  BUFx4f_ASAP7_75t_R register___U3006 ( .A(register__n11843), .Y(register__n11839) );
  HB1xp67_ASAP7_75t_R register___U3007 ( .A(register__n12528), .Y(register__n5748) );
  INVx1_ASAP7_75t_R register___U3008 ( .A(register__n12677), .Y(register__n6994) );
  BUFx6f_ASAP7_75t_R register___U3009 ( .A(register__net141997), .Y(register__net63352) );
  INVxp67_ASAP7_75t_R register___U3010 ( .A(register__net63362), .Y(register__net63330) );
  INVx1_ASAP7_75t_R register___U3011 ( .A(register__net63382), .Y(register__net63346) );
  INVx4_ASAP7_75t_R register___U3012 ( .A(register__net63334), .Y(register__net100610) );
  HB1xp67_ASAP7_75t_R register___U3013 ( .A(register__n4207), .Y(register__n4206) );
  HB1xp67_ASAP7_75t_R register___U3014 ( .A(register__n5766), .Y(register__n5765) );
  INVx1_ASAP7_75t_R register___U3015 ( .A(register__n1792), .Y(register__n1618) );
  BUFx4f_ASAP7_75t_R register___U3016 ( .A(register__net64038), .Y(register__net64040) );
  NOR2xp67_ASAP7_75t_R register___U3017 ( .A(register__n2770), .B(register__n2771), .Y(register__n13194) );
  BUFx12f_ASAP7_75t_R register___U3018 ( .A(register__n3993), .Y(register__n12044) );
  AO22x2_ASAP7_75t_R register___U3019 ( .A1(register__net64972), .A2(register__n1618), .B1(register__n846), .B2(register__n1647), 
        .Y(register__n845) );
  CKINVDCx20_ASAP7_75t_R register___U3020 ( .A(register__n9923), .Y(register__n846) );
  CKINVDCx5p33_ASAP7_75t_R register___U3021 ( .A(register__net64972), .Y(register__net64938) );
  AO22x1_ASAP7_75t_R register___U3022 ( .A1(register__n9816), .A2(register__C6422_net70498), .B1(register__n10227), 
        .B2(register__net126625), .Y(register__n10753) );
  NAND2xp33_ASAP7_75t_R register___U3023 ( .A(register__net89909), .B(register__net126625), .Y(register__n2366) );
  AO22x1_ASAP7_75t_R register___U3024 ( .A1(register__n9579), .A2(register__n1771), .B1(register__n9999), .B2(register__net126625), .Y(register__n10971) );
  AO22x1_ASAP7_75t_R register___U3025 ( .A1(register__n8347), .A2(register__net121619), .B1(register__n8803), .B2(
        net126625), .Y(register__n10857) );
  AO22x1_ASAP7_75t_R register___U3026 ( .A1(register__n9828), .A2(register__net121619), .B1(register__n10243), .B2(
        net126625), .Y(register__n10904) );
  AO22x1_ASAP7_75t_R register___U3027 ( .A1(register__n9855), .A2(register__n1771), .B1(register__n10281), .B2(
        C6422_net70534), .Y(register__n11032) );
  AO22x1_ASAP7_75t_R register___U3028 ( .A1(register__n7400), .A2(register__net121619), .B1(register__n5648), .B2(
        net126625), .Y(register__n10948) );
  AO22x1_ASAP7_75t_R register___U3029 ( .A1(register__net90213), .A2(register__n1771), .B1(register__net89565), .B2(
        net126625), .Y(register__n11095) );
  AO22x1_ASAP7_75t_R register___U3030 ( .A1(register__n9836), .A2(register__net121619), .B1(register__n10253), .B2(
        net126625), .Y(register__n10992) );
  AO22x1_ASAP7_75t_R register___U3031 ( .A1(register__n10519), .A2(register__net121619), .B1(register__n5206), .B2(
        net126625), .Y(register__n10881) );
  INVx1_ASAP7_75t_R register___U3032 ( .A(register__n12719), .Y(register__n847) );
  INVx1_ASAP7_75t_R register___U3033 ( .A(register__n1787), .Y(register__n1636) );
  AO22x1_ASAP7_75t_R register___U3034 ( .A1(register__net64056), .A2(register__n11802), .B1(register__n2705), .B2(register__n109), 
        .Y(register__n1606) );
  INVxp33_ASAP7_75t_R register___U3035 ( .A(register__n1645), .Y(register__n11811) );
  INVxp33_ASAP7_75t_R register___U3036 ( .A(register__n1792), .Y(register__n1621) );
  INVxp33_ASAP7_75t_R register___U3037 ( .A(register__n3832), .Y(register__n1779) );
  INVxp33_ASAP7_75t_R register___U3038 ( .A(register__n3832), .Y(register__n1630) );
  INVxp67_ASAP7_75t_R register___U3039 ( .A(register__n11811), .Y(register__n11893) );
  HB1xp67_ASAP7_75t_R register___U3040 ( .A(register__n11077), .Y(register__n4995) );
  AO22x1_ASAP7_75t_R register___U3041 ( .A1(register__n3), .A2(register__n10505), .B1(register__n10425), .B2(register__n1578), 
        .Y(register__n11077) );
  HB1xp67_ASAP7_75t_R register___U3042 ( .A(register__n13214), .Y(register__n3894) );
  INVxp67_ASAP7_75t_R register___U3043 ( .A(register__n13168), .Y(register__n848) );
  HB1xp67_ASAP7_75t_R register___U3044 ( .A(register__n12938), .Y(register__n3743) );
  HB1xp67_ASAP7_75t_R register___U3045 ( .A(register__n3656), .Y(register__n3655) );
  INVx4_ASAP7_75t_R register___U3046 ( .A(register__n3669), .Y(register__n11922) );
  HB1xp67_ASAP7_75t_R register___U3047 ( .A(register__n13318), .Y(register__n4061) );
  INVxp33_ASAP7_75t_R register___U3048 ( .A(register__n10518), .Y(register__n1947) );
  INVx1_ASAP7_75t_R register___U3049 ( .A(register__n11329), .Y(register__n8278) );
  INVx2_ASAP7_75t_R register___U3050 ( .A(register__n8278), .Y(register__n1178) );
  HB1xp67_ASAP7_75t_R register___U3051 ( .A(register__net122862), .Y(register__net125804) );
  INVx1_ASAP7_75t_R register___U3052 ( .A(register__n13263), .Y(register__n850) );
  BUFx6f_ASAP7_75t_R register___U3053 ( .A(register__n11750), .Y(register__n3295) );
  BUFx12f_ASAP7_75t_R register___U3054 ( .A(register__n3260), .Y(register__n3503) );
  INVx1_ASAP7_75t_R register___U3055 ( .A(register__n12701), .Y(register__n851) );
  INVx1_ASAP7_75t_R register___U3056 ( .A(register__n12797), .Y(register__n852) );
  INVx1_ASAP7_75t_R register___U3057 ( .A(register__n13077), .Y(register__n853) );
  INVx1_ASAP7_75t_R register___U3058 ( .A(register__n12704), .Y(register__n854) );
  INVx3_ASAP7_75t_R register___U3059 ( .A(register__n12061), .Y(register__n855) );
  INVx2_ASAP7_75t_R register___U3060 ( .A(register__n12075), .Y(register__n12061) );
  INVxp33_ASAP7_75t_R register___U3061 ( .A(register__n1080), .Y(register__n11716) );
  AOI22xp33_ASAP7_75t_R register___U3062 ( .A1(register__n9891), .A2(register__C6423_net61340), .B1(register__n9321), 
        .B2(register__C6423_net69198), .Y(register__n1080) );
  INVx2_ASAP7_75t_R register___U3063 ( .A(register__net93286), .Y(register__net122602) );
  BUFx2_ASAP7_75t_R register___U3064 ( .A(register__net122603), .Y(register__net93286) );
  HB1xp67_ASAP7_75t_R register___U3065 ( .A(register__C6423_net60474), .Y(register__net122603) );
  BUFx12f_ASAP7_75t_R register___U3066 ( .A(register__n11752), .Y(register__n3277) );
  NOR2xp33_ASAP7_75t_R register___U3067 ( .A(register__n1995), .B(register__C6422_net59704), .Y(register__n857) );
  AND2x2_ASAP7_75t_R register___U3068 ( .A(register__n11260), .B(register__n11262), .Y(register__n859) );
  AND3x1_ASAP7_75t_R register___U3069 ( .A(register__n11261), .B(register__n859), .C(register__n493), .Y(register__n8643) );
  INVx2_ASAP7_75t_R register___U3070 ( .A(register__net88949), .Y(register__C6422_net59703) );
  INVx3_ASAP7_75t_R register___U3071 ( .A(register__net91523), .Y(register__C6422_net59704) );
  HB1xp67_ASAP7_75t_R register___U3072 ( .A(register__C6423_net60623), .Y(register__net113304) );
  AND3x2_ASAP7_75t_R register___U3073 ( .A(register__n1329), .B(register__n7053), .C(register__n1328), .Y(register__n11262) );
  INVx1_ASAP7_75t_R register___U3074 ( .A(register__n1974), .Y(register__n2892) );
  BUFx12f_ASAP7_75t_R register___U3075 ( .A(register__n11787), .Y(register__n2891) );
  AND2x2_ASAP7_75t_R register___U3076 ( .A(register__n10884), .B(register__n10885), .Y(register__n860) );
  AND3x1_ASAP7_75t_R register___U3077 ( .A(register__n860), .B(register__n8291), .C(register__n10883), .Y(register__n7940) );
  INVxp67_ASAP7_75t_R register___U3078 ( .A(register__n10886), .Y(register__n8291) );
  BUFx12f_ASAP7_75t_R register___U3079 ( .A(register__n8561), .Y(register__n12074) );
  BUFx12f_ASAP7_75t_R register___U3080 ( .A(register__n855), .Y(register__n12071) );
  INVx1_ASAP7_75t_R register___U3081 ( .A(register__net64886), .Y(register__net64852) );
  NOR2x2_ASAP7_75t_R register___U3082 ( .A(register__n12058), .B(register__n2812), .Y(register__n2795) );
  NOR2x1p5_ASAP7_75t_R register___U3083 ( .A(register__n2795), .B(register__n73), .Y(register__n12879) );
  NAND2x1p5_ASAP7_75t_R register___U3084 ( .A(register__n862), .B(register__n863), .Y(register__n1007) );
  HB1xp67_ASAP7_75t_R register___U3085 ( .A(register__n10515), .Y(register__n6605) );
  HB1xp67_ASAP7_75t_R register___U3086 ( .A(register__n10513), .Y(register__n8202) );
  BUFx3_ASAP7_75t_R register___U3087 ( .A(register__n5337), .Y(register__n5336) );
  AND2x2_ASAP7_75t_R register___U3088 ( .A(register__n9182), .B(register__n864), .Y(register__n10657) );
  INVx1_ASAP7_75t_R register___U3089 ( .A(register__n10666), .Y(register__n9182) );
  BUFx6f_ASAP7_75t_R register___U3090 ( .A(register__n3647), .Y(register__n8245) );
  INVx2_ASAP7_75t_R register___U3091 ( .A(register__n12271), .Y(register__n12258) );
  BUFx6f_ASAP7_75t_R register___U3092 ( .A(register__n8245), .Y(register__n12271) );
  NOR2x1p5_ASAP7_75t_R register___U3093 ( .A(register__net98142), .B(register__net107120), .Y(register__n2426) );
  HB1xp67_ASAP7_75t_R register___U3094 ( .A(register__n13046), .Y(register__n5080) );
  HB1xp67_ASAP7_75t_R register___U3095 ( .A(register__n5760), .Y(register__n5759) );
  INVx1_ASAP7_75t_R register___U3096 ( .A(register__n12549), .Y(register__n865) );
  INVx1_ASAP7_75t_R register___U3097 ( .A(register__n10614), .Y(register__n866) );
  BUFx3_ASAP7_75t_R register___U3098 ( .A(register__n11241), .Y(register__n5995) );
  BUFx12f_ASAP7_75t_R register___U3099 ( .A(register__n8563), .Y(register__n12073) );
  BUFx4f_ASAP7_75t_R register___U3100 ( .A(register__net102927), .Y(register__net64890) );
  OR2x2_ASAP7_75t_R register___U3101 ( .A(register__n1903), .B(register__n2703), .Y(register__n867) );
  NOR2xp33_ASAP7_75t_R register___U3102 ( .A(register__n2710), .B(register__n2713), .Y(register__n868) );
  NOR3xp33_ASAP7_75t_R register___U3103 ( .A(register__n869), .B(register__n2706), .C(register__n2709), .Y(register__n2732) );
  INVxp67_ASAP7_75t_R register___U3104 ( .A(register__n868), .Y(register__n869) );
  INVxp33_ASAP7_75t_R register___U3105 ( .A(register__net89389), .Y(register__n2703) );
  NOR2xp33_ASAP7_75t_R register___U3106 ( .A(register__n2708), .B(register__n_cell_125074_net170535), .Y(
        n2710) );
  NOR2xp33_ASAP7_75t_R register___U3107 ( .A(register__n2711), .B(register__n276), .Y(register__n2713) );
  INVx1_ASAP7_75t_R register___U3108 ( .A(register__n13224), .Y(register__n870) );
  BUFx6f_ASAP7_75t_R register___U3109 ( .A(register__n11733), .Y(register__n11852) );
  INVx6_ASAP7_75t_R register___U3110 ( .A(register__net64418), .Y(register__net127722) );
  INVx1_ASAP7_75t_R register___U3111 ( .A(register__n2016), .Y(register__n2018) );
  INVx1_ASAP7_75t_R register___U3112 ( .A(register__n2018), .Y(register__n1915) );
  BUFx4f_ASAP7_75t_R register___U3113 ( .A(register__n3475), .Y(register__n12477) );
  BUFx3_ASAP7_75t_R register___U3114 ( .A(register__n3392), .Y(register__n3267) );
  BUFx12f_ASAP7_75t_R register___U3115 ( .A(register__n3191), .Y(register__n11734) );
  INVxp67_ASAP7_75t_R register___U3116 ( .A(register__n2931), .Y(register__n4048) );
  HB1xp67_ASAP7_75t_R register___U3117 ( .A(register__n12903), .Y(register__n2931) );
  INVx6_ASAP7_75t_R register___U3118 ( .A(register__n4836), .Y(register__n12323) );
  AOI21xp33_ASAP7_75t_R register___U3119 ( .A1(register__net88817), .A2(register__net109611), .B(register__n2510), .Y(
        n2512) );
  AOI21xp33_ASAP7_75t_R register___U3120 ( .A1(register__net88857), .A2(register__C6423_net60464), .B(register__n2691), 
        .Y(register__n2719) );
  AO22x1_ASAP7_75t_R register___U3121 ( .A1(register__n10434), .A2(register__n883), .B1(register__n10421), .B2(
        net122862), .Y(register__n11357) );
  INVxp67_ASAP7_75t_R register___U3122 ( .A(register__n1767), .Y(register__n1302) );
  INVxp67_ASAP7_75t_R register___U3123 ( .A(register__n4086), .Y(register__n4990) );
  BUFx12f_ASAP7_75t_R register___U3124 ( .A(register__n3947), .Y(register__n5929) );
  INVx4_ASAP7_75t_R register___U3125 ( .A(register__n1403), .Y(register__n3947) );
  NAND3x1_ASAP7_75t_R register___U3126 ( .A(register__n1297), .B(register__n10840), .C(register__n5915), .Y(register__n872) );
  AND3x2_ASAP7_75t_R register___U3127 ( .A(register__n11143), .B(register__n11132), .C(IF_ID_rs1[2]), 
        .Y(register__n11131) );
  HB1xp67_ASAP7_75t_R register___U3128 ( .A(register__n12162), .Y(register__n4849) );
  BUFx4f_ASAP7_75t_R register___U3129 ( .A(register__n112), .Y(register__net99872) );
  BUFx12f_ASAP7_75t_R register___U3130 ( .A(write_data[15]), .Y(register__net64062) );
  HB1xp67_ASAP7_75t_R register___U3131 ( .A(register__n13218), .Y(register__n4516) );
  HB1xp67_ASAP7_75t_R register___U3132 ( .A(register__n12706), .Y(register__n3687) );
  INVx1_ASAP7_75t_R register___U3133 ( .A(register__n12565), .Y(register__n873) );
  HB1xp67_ASAP7_75t_R register___U3134 ( .A(register__n12191), .Y(register__n12179) );
  HB1xp67_ASAP7_75t_R register___U3135 ( .A(register__n12191), .Y(register__n12184) );
  HB1xp67_ASAP7_75t_R register___U3136 ( .A(register__n12191), .Y(register__n12183) );
  INVx1_ASAP7_75t_R register___U3137 ( .A(register__n12184), .Y(register__n12172) );
  INVxp67_ASAP7_75t_R register___U3138 ( .A(register__n12183), .Y(register__n12167) );
  HB1xp67_ASAP7_75t_R register___U3139 ( .A(register__n12735), .Y(register__n3782) );
  BUFx6f_ASAP7_75t_R register___U3140 ( .A(register__n3917), .Y(register__n3877) );
  BUFx3_ASAP7_75t_R register___U3141 ( .A(register__n12022), .Y(register__n3073) );
  INVx1_ASAP7_75t_R register___U3142 ( .A(register__n3073), .Y(register__n1025) );
  INVxp67_ASAP7_75t_R register___U3143 ( .A(register__n1915), .Y(register__n1916) );
  INVxp67_ASAP7_75t_R register___U3144 ( .A(register__n1915), .Y(register__n1917) );
  AOI22xp33_ASAP7_75t_R register___U3145 ( .A1(register__n12362), .A2(register__n2135), .B1(register__n874), .B2(register__n1576), 
        .Y(register__n12898) );
  CKINVDCx20_ASAP7_75t_R register___U3146 ( .A(register__n8817), .Y(register__n874) );
  INVx2_ASAP7_75t_R register___U3147 ( .A(register__n12357), .Y(register__n12344) );
  BUFx3_ASAP7_75t_R register___U3148 ( .A(register__n5348), .Y(register__n12362) );
  BUFx12f_ASAP7_75t_R register___U3149 ( .A(register__n3336), .Y(register__n3335) );
  HB1xp67_ASAP7_75t_R register___U3150 ( .A(register__n2984), .Y(register__n2968) );
  NAND2xp5_ASAP7_75t_R register___U3151 ( .A(register__n12034), .B(register__n2968), .Y(register__n1956) );
  HB1xp67_ASAP7_75t_R register___U3152 ( .A(register__n4745), .Y(register__n12295) );
  AND3x2_ASAP7_75t_R register___U3153 ( .A(register__n2233), .B(register__n5441), .C(register__n11721), .Y(register__n877) );
  OAI22xp33_ASAP7_75t_R register___U3154 ( .A1(register__n12377), .A2(register__n7327), .B1(register__n9579), .B2(register__n5929), .Y(register__n878) );
  AO22x1_ASAP7_75t_R register___U3155 ( .A1(register__n10440), .A2(register__n3), .B1(register__n10469), .B2(register__n281), .Y(
        n10905) );
  CKINVDCx20_ASAP7_75t_R register___U3156 ( .A(register__n120), .Y(register__n879) );
  OR2x2_ASAP7_75t_R register___U3157 ( .A(register__n2659), .B(register__n367), .Y(register__n881) );
  NAND2xp33_ASAP7_75t_R register___U3158 ( .A(register__n881), .B(register__n2683), .Y(register__n2684) );
  INVxp33_ASAP7_75t_R register___U3159 ( .A(register__net89413), .Y(register__n2659) );
  AOI211x1_ASAP7_75t_R register___U3160 ( .A1(register__net90877), .A2(register__C6423_net72255), .B(register__n2443), 
        .C(register__n2439), .Y(register__n2442) );
  BUFx3_ASAP7_75t_R register___U3161 ( .A(register__net125426), .Y(register__net138603) );
  BUFx4f_ASAP7_75t_R register___U3162 ( .A(register__net122599), .Y(register__net137440) );
  BUFx3_ASAP7_75t_R register___U3163 ( .A(register__net137440), .Y(register__net93282) );
  INVx1_ASAP7_75t_R register___U3164 ( .A(register__C6423_net72243), .Y(register__C6423_net72255) );
  BUFx2_ASAP7_75t_R register___U3165 ( .A(register__net137440), .Y(register__net139572) );
  BUFx6f_ASAP7_75t_R register___U3166 ( .A(register__net93282), .Y(register__net128003) );
  BUFx6f_ASAP7_75t_R register___U3167 ( .A(register__net139047), .Y(register__net125425) );
  INVx2_ASAP7_75t_R register___U3168 ( .A(register__net125425), .Y(register__C6423_net72245) );
  INVx4_ASAP7_75t_R register___U3169 ( .A(register__net136856), .Y(register__C6423_net72242) );
  HB1xp67_ASAP7_75t_R register___U3170 ( .A(register__n5034), .Y(register__n4283) );
  HB1xp67_ASAP7_75t_R register___U3171 ( .A(register__n5034), .Y(register__n12102) );
  HB1xp67_ASAP7_75t_R register___U3172 ( .A(register__n5034), .Y(register__n12106) );
  HB1xp67_ASAP7_75t_R register___U3173 ( .A(register__n5034), .Y(register__n12101) );
  AOI22x1_ASAP7_75t_R register___U3174 ( .A1(register__net64886), .A2(register__n534), .B1(register__n1097), .B2(register__n1098), 
        .Y(register__n12795) );
  CKINVDCx10_ASAP7_75t_R register___U3175 ( .A(register__n3737), .Y(register__n3735) );
  BUFx12f_ASAP7_75t_R register___U3176 ( .A(register__n3360), .Y(register__n3737) );
  INVx1_ASAP7_75t_R register___U3177 ( .A(register__n12594), .Y(register__n886) );
  BUFx3_ASAP7_75t_R register___U3178 ( .A(register__n11125), .Y(register__n5156) );
  HB1xp67_ASAP7_75t_R register___U3179 ( .A(register__n4087), .Y(register__n4086) );
  INVxp67_ASAP7_75t_R register___U3180 ( .A(register__n1268), .Y(register__n12762) );
  AO22x1_ASAP7_75t_R register___U3181 ( .A1(register__net64048), .A2(register__n1620), .B1(register__n1269), .B2(register__n1643), 
        .Y(register__n1268) );
  BUFx12f_ASAP7_75t_R register___U3182 ( .A(register__n11764), .Y(register__n887) );
  BUFx6f_ASAP7_75t_R register___U3183 ( .A(register__n11764), .Y(register__n888) );
  INVx2_ASAP7_75t_R register___U3184 ( .A(register__n4968), .Y(register__n891) );
  INVx2_ASAP7_75t_R register___U3185 ( .A(register__n4968), .Y(register__n892) );
  INVx6_ASAP7_75t_R register___U3186 ( .A(register__n887), .Y(register__n896) );
  INVx2_ASAP7_75t_R register___U3187 ( .A(register__n887), .Y(register__n897) );
  INVx2_ASAP7_75t_R register___U3188 ( .A(register__n887), .Y(register__n898) );
  INVx2_ASAP7_75t_R register___U3189 ( .A(register__n887), .Y(register__n899) );
  INVx2_ASAP7_75t_R register___U3190 ( .A(register__n887), .Y(register__n900) );
  INVx2_ASAP7_75t_R register___U3191 ( .A(register__n888), .Y(register__n902) );
  INVx2_ASAP7_75t_R register___U3192 ( .A(register__n888), .Y(register__n903) );
  INVx2_ASAP7_75t_R register___U3193 ( .A(register__n888), .Y(register__n904) );
  INVx2_ASAP7_75t_R register___U3194 ( .A(register__n888), .Y(register__n905) );
  INVx2_ASAP7_75t_R register___U3195 ( .A(register__n888), .Y(register__n906) );
  INVx2_ASAP7_75t_R register___U3196 ( .A(register__n888), .Y(register__n907) );
  NAND2xp67_ASAP7_75t_R register___U3197 ( .A(register__n910), .B(register__n909), .Y(read_reg_data_2[24]) );
  CKINVDCx20_ASAP7_75t_R register___U3198 ( .A(register__n1251), .Y(register__n909) );
  INVxp33_ASAP7_75t_R register___U3199 ( .A(register__net122579), .Y(register__n918) );
  INVxp67_ASAP7_75t_R register___U3200 ( .A(register__n913), .Y(register__n924) );
  INVxp33_ASAP7_75t_R register___U3201 ( .A(register__n918), .Y(register__n933) );
  INVxp33_ASAP7_75t_R register___U3202 ( .A(register__n918), .Y(register__n934) );
  HB1xp67_ASAP7_75t_R register___U3203 ( .A(register__net122579), .Y(register__net118097) );
  HB1xp67_ASAP7_75t_R register___U3204 ( .A(register__net118097), .Y(register__net128096) );
  BUFx12f_ASAP7_75t_R register___U3205 ( .A(register__n2970), .Y(register__n2965) );
  INVx1_ASAP7_75t_R register___U3206 ( .A(register__n12509), .Y(register__n2246) );
  AO22x1_ASAP7_75t_R register___U3207 ( .A1(register__n9728), .A2(register__net109849), .B1(register__n10183), .B2(register__n634), .Y(register__n11319) );
  INVxp33_ASAP7_75t_R register___U3208 ( .A(register__n4950), .Y(register__n8702) );
  INVx1_ASAP7_75t_R register___U3209 ( .A(register__n4371), .Y(register__n7596) );
  AND2x2_ASAP7_75t_R register___U3210 ( .A(register__n4003), .B(register__n7931), .Y(register__n935) );
  AND2x2_ASAP7_75t_R register___U3211 ( .A(register__n1229), .B(register__n935), .Y(register__n11343) );
  INVxp67_ASAP7_75t_R register___U3212 ( .A(register__n2965), .Y(register__n1599) );
  BUFx6f_ASAP7_75t_R register___U3213 ( .A(register__n3425), .Y(register__n3449) );
  AO22x1_ASAP7_75t_R register___U3214 ( .A1(register__n9849), .A2(register__C6423_net61333), .B1(register__n8523), .B2(
        C6423_net61331), .Y(register__n11361) );
  HB1xp67_ASAP7_75t_R register___U3215 ( .A(register__n11361), .Y(register__n4557) );
  OAI22xp33_ASAP7_75t_R register___U3216 ( .A1(register__net62984), .A2(register__n1988), .B1(register__n8353), .B2(
        n2984), .Y(register__n936) );
  INVx1_ASAP7_75t_R register___U3217 ( .A(register__n12723), .Y(register__n937) );
  BUFx2_ASAP7_75t_R register___U3218 ( .A(register__n4372), .Y(register__n4371) );
  INVxp67_ASAP7_75t_R register___U3219 ( .A(register__n13105), .Y(register__n5902) );
  INVx1_ASAP7_75t_R register___U3220 ( .A(register__n12640), .Y(register__n938) );
  INVxp67_ASAP7_75t_R register___U3221 ( .A(register__n4677), .Y(register__n8615) );
  HB1xp67_ASAP7_75t_R register___U3222 ( .A(register__n12899), .Y(register__n2920) );
  BUFx3_ASAP7_75t_R register___U3223 ( .A(register__n4953), .Y(register__n3392) );
  AOI22xp33_ASAP7_75t_R register___U3224 ( .A1(register__n12387), .A2(register__n1734), .B1(register__n939), .B2(register__n1724), 
        .Y(register__n13247) );
  CKINVDCx20_ASAP7_75t_R register___U3225 ( .A(register__n9999), .Y(register__n939) );
  BUFx2_ASAP7_75t_R register___U3226 ( .A(register__n4954), .Y(register__n4953) );
  NOR2xp33_ASAP7_75t_R register___U3227 ( .A(register__n2080), .B(register__n6217), .Y(register__n940) );
  NOR2xp33_ASAP7_75t_R register___U3228 ( .A(register__n11247), .B(register__net112580), .Y(register__n942) );
  NOR3xp33_ASAP7_75t_R register___U3229 ( .A(register__n940), .B(register__n941), .C(register__n942), .Y(register__n10615) );
  HB1xp67_ASAP7_75t_R register___U3230 ( .A(register__n10621), .Y(register__n6217) );
  HB1xp67_ASAP7_75t_R register___U3231 ( .A(register__n5626), .Y(register__n5625) );
  BUFx3_ASAP7_75t_R register___U3232 ( .A(register__net138603), .Y(register__net139047) );
  OAI21xp33_ASAP7_75t_R register___U3233 ( .A1(register__n488), .A2(register__n2432), .B(register__n2453), .Y(register__n2452) );
  AO22x1_ASAP7_75t_R register___U3234 ( .A1(register__n9730), .A2(register__n481), .B1(register__n10098), .B2(register__n635), 
        .Y(register__n11364) );
  AO22x1_ASAP7_75t_R register___U3235 ( .A1(register__n9646), .A2(register__net109849), .B1(register__n9973), .B2(register__n640), 
        .Y(register__n11493) );
  AO22x1_ASAP7_75t_R register___U3236 ( .A1(register__net90901), .A2(register__n482), .B1(register__net89993), .B2(
        C6423_net61348), .Y(register__n11277) );
  INVx1_ASAP7_75t_R register___U3237 ( .A(register__n12753), .Y(register__n943) );
  INVx6_ASAP7_75t_R register___U3238 ( .A(register__n11825), .Y(register__n11907) );
  INVx3_ASAP7_75t_R register___U3239 ( .A(register__n2285), .Y(register__n11827) );
  HB1xp67_ASAP7_75t_R register___U3240 ( .A(register__n13057), .Y(register__n5756) );
  INVx1_ASAP7_75t_R register___U3241 ( .A(register__n13176), .Y(register__n944) );
  AOI22xp33_ASAP7_75t_R register___U3242 ( .A1(register__C6422_net59538), .A2(register__n9541), .B1(
        C6422_net59540), .B2(register__n7395), .Y(register__n10785) );
  INVx1_ASAP7_75t_R register___U3243 ( .A(register__n13162), .Y(register__n945) );
  BUFx6f_ASAP7_75t_R register___U3244 ( .A(register__n11843), .Y(register__n3359) );
  BUFx12f_ASAP7_75t_R register___U3245 ( .A(register__n12048), .Y(register__n3993) );
  HB1xp67_ASAP7_75t_R register___U3246 ( .A(register__n4678), .Y(register__n4677) );
  INVx1_ASAP7_75t_R register___U3247 ( .A(register__n12552), .Y(register__n947) );
  INVx1_ASAP7_75t_R register___U3248 ( .A(register__n13151), .Y(register__n948) );
  INVx1_ASAP7_75t_R register___U3249 ( .A(register__n13157), .Y(register__n949) );
  INVx1_ASAP7_75t_R register___U3250 ( .A(register__n13152), .Y(register__n950) );
  BUFx12f_ASAP7_75t_R register___U3251 ( .A(register__C6423_net60464), .Y(register__net109611) );
  AOI21xp33_ASAP7_75t_R register___U3252 ( .A1(register__C6423_net60464), .A2(register__net88957), .B(register__n2424), 
        .Y(register__n2444) );
  BUFx12f_ASAP7_75t_R register___U3253 ( .A(register__n3543), .Y(register__n4633) );
  CKINVDCx10_ASAP7_75t_R register___U3254 ( .A(register__n12126), .Y(register__n12125) );
  HB1xp67_ASAP7_75t_R register___U3255 ( .A(register__n12126), .Y(register__n12132) );
  INVx1_ASAP7_75t_R register___U3256 ( .A(register__n3944), .Y(register__n955) );
  INVx1_ASAP7_75t_R register___U3257 ( .A(register__n3944), .Y(register__n956) );
  INVx6_ASAP7_75t_R register___U3258 ( .A(register__n11765), .Y(register__n958) );
  CKINVDCx5p33_ASAP7_75t_R register___U3259 ( .A(register__n11765), .Y(register__n959) );
  INVx5_ASAP7_75t_R register___U3260 ( .A(register__n11765), .Y(register__n960) );
  INVx1_ASAP7_75t_R register___U3261 ( .A(register__n13011), .Y(register__n961) );
  CKINVDCx5p33_ASAP7_75t_R register___U3262 ( .A(register__n3944), .Y(register__n11765) );
  INVx1_ASAP7_75t_R register___U3263 ( .A(register__n13149), .Y(register__n962) );
  INVx1_ASAP7_75t_R register___U3264 ( .A(register__n13160), .Y(register__n963) );
  INVx1_ASAP7_75t_R register___U3265 ( .A(register__n13175), .Y(register__n964) );
  INVx2_ASAP7_75t_R register___U3266 ( .A(register__n4001), .Y(register__n12114) );
  BUFx12f_ASAP7_75t_R register___U3267 ( .A(register__n3839), .Y(register__n4001) );
  NOR2xp33_ASAP7_75t_R register___U3268 ( .A(register__net62656), .B(register__n103), .Y(register__n965) );
  NOR2xp33_ASAP7_75t_R register___U3269 ( .A(register__n7723), .B(register__n1151), .Y(register__n966) );
  NOR2xp33_ASAP7_75t_R register___U3270 ( .A(register__n965), .B(register__n966), .Y(register__n13148) );
  INVxp67_ASAP7_75t_R register___U3271 ( .A(register__n13148), .Y(register__n967) );
  INVx1_ASAP7_75t_R register___U3272 ( .A(register__n13171), .Y(register__n968) );
  INVx1_ASAP7_75t_R register___U3273 ( .A(register__n7633), .Y(register__n969) );
  INVx1_ASAP7_75t_R register___U3274 ( .A(register__n7633), .Y(register__n970) );
  INVx1_ASAP7_75t_R register___U3275 ( .A(register__n7633), .Y(register__n971) );
  INVx1_ASAP7_75t_R register___U3276 ( .A(register__n7633), .Y(register__n972) );
  INVxp67_ASAP7_75t_R register___U3277 ( .A(register__n7633), .Y(register__n973) );
  INVxp67_ASAP7_75t_R register___U3278 ( .A(register__n7633), .Y(register__n974) );
  INVxp67_ASAP7_75t_R register___U3279 ( .A(register__n7633), .Y(register__n975) );
  INVxp67_ASAP7_75t_R register___U3280 ( .A(register__n1812), .Y(register__n977) );
  INVx1_ASAP7_75t_R register___U3281 ( .A(register__n1811), .Y(register__n978) );
  INVxp33_ASAP7_75t_R register___U3282 ( .A(register__n1808), .Y(register__n979) );
  INVxp33_ASAP7_75t_R register___U3283 ( .A(register__n1807), .Y(register__n980) );
  INVxp33_ASAP7_75t_R register___U3284 ( .A(register__n1809), .Y(register__n981) );
  INVxp67_ASAP7_75t_R register___U3285 ( .A(register__n1810), .Y(register__n982) );
  INVxp33_ASAP7_75t_R register___U3286 ( .A(register__n1814), .Y(register__n983) );
  INVx1_ASAP7_75t_R register___U3287 ( .A(register__n3711), .Y(register__n985) );
  INVxp67_ASAP7_75t_R register___U3288 ( .A(register__n1818), .Y(register__n986) );
  INVx1_ASAP7_75t_R register___U3289 ( .A(register__n3709), .Y(register__n988) );
  INVxp67_ASAP7_75t_R register___U3290 ( .A(register__n1820), .Y(register__n991) );
  INVxp67_ASAP7_75t_R register___U3291 ( .A(register__n1822), .Y(register__n992) );
  INVxp67_ASAP7_75t_R register___U3292 ( .A(register__n4955), .Y(register__n993) );
  INVx2_ASAP7_75t_R register___U3293 ( .A(register__n11875), .Y(register__n994) );
  INVxp67_ASAP7_75t_R register___U3294 ( .A(register__n1824), .Y(register__n995) );
  INVxp67_ASAP7_75t_R register___U3295 ( .A(register__n1826), .Y(register__n996) );
  INVx2_ASAP7_75t_R register___U3296 ( .A(register__n3168), .Y(register__n997) );
  INVx2_ASAP7_75t_R register___U3297 ( .A(register__n3169), .Y(register__n998) );
  INVxp67_ASAP7_75t_R register___U3298 ( .A(register__n1830), .Y(register__n999) );
  INVx2_ASAP7_75t_R register___U3299 ( .A(register__n11874), .Y(register__n1000) );
  INVxp67_ASAP7_75t_R register___U3300 ( .A(register__n1828), .Y(register__n1001) );
  INVx1_ASAP7_75t_R register___U3301 ( .A(register__n4840), .Y(register__n1002) );
  INVx1_ASAP7_75t_R register___U3302 ( .A(register__n1832), .Y(register__n1003) );
  INVx6_ASAP7_75t_R register___U3303 ( .A(register__n5355), .Y(register__n1004) );
  INVx1_ASAP7_75t_R register___U3304 ( .A(register__n1834), .Y(register__n1005) );
  CKINVDCx10_ASAP7_75t_R register___U3305 ( .A(register__n5515), .Y(register__n5516) );
  INVxp67_ASAP7_75t_R register___U3306 ( .A(register__n1815), .Y(register__n1816) );
  INVxp33_ASAP7_75t_R register___U3307 ( .A(register__n1819), .Y(register__n1820) );
  INVxp33_ASAP7_75t_R register___U3308 ( .A(register__n1821), .Y(register__n1822) );
  INVxp33_ASAP7_75t_R register___U3309 ( .A(register__n1823), .Y(register__n1824) );
  BUFx12f_ASAP7_75t_R register___U3310 ( .A(register__n9379), .Y(register__n3168) );
  HB1xp67_ASAP7_75t_R register___U3311 ( .A(register__n9379), .Y(register__n3169) );
  INVxp33_ASAP7_75t_R register___U3312 ( .A(register__n1827), .Y(register__n1828) );
  HB1xp67_ASAP7_75t_R register___U3313 ( .A(register__n11875), .Y(register__n4840) );
  INVxp67_ASAP7_75t_R register___U3314 ( .A(register__n11875), .Y(register__n1827) );
  INVxp33_ASAP7_75t_R register___U3315 ( .A(register__n4955), .Y(register__n1829) );
  INVxp67_ASAP7_75t_R register___U3316 ( .A(register__n9379), .Y(register__n1825) );
  INVx2_ASAP7_75t_R register___U3317 ( .A(register__n11874), .Y(register__n1833) );
  INVx6_ASAP7_75t_R register___U3318 ( .A(register__n12073), .Y(register__n12060) );
  INVx1_ASAP7_75t_R register___U3319 ( .A(register__n12879), .Y(register__n2272) );
  HB1xp67_ASAP7_75t_R register___U3320 ( .A(register__n12049), .Y(register__n12045) );
  NOR4xp75_ASAP7_75t_R register___U3321 ( .A(register__n1007), .B(register__n11044), .C(register__n3617), .D(register__n11046), 
        .Y(register__n11036) );
  INVx4_ASAP7_75t_R register___U3322 ( .A(register__net97185), .Y(register__net105518) );
  INVx1_ASAP7_75t_R register___U3323 ( .A(register__n13155), .Y(register__n1009) );
  AO22x1_ASAP7_75t_R register___U3324 ( .A1(register__n9613), .A2(register__C6423_net61343), .B1(register__n10080), 
        .B2(register__net129787), .Y(register__n11486) );
  AO22x1_ASAP7_75t_R register___U3325 ( .A1(register__n8757), .A2(register__C6423_net61343), .B1(register__n8084), .B2(
        C6423_net69274), .Y(register__n11252) );
  AO22x1_ASAP7_75t_R register___U3326 ( .A1(register__n9615), .A2(register__C6423_net61343), .B1(register__n10084), 
        .B2(register__net129787), .Y(register__n11232) );
  AO22x1_ASAP7_75t_R register___U3327 ( .A1(register__n8809), .A2(register__C6423_net61343), .B1(register__n8353), .B2(
        net129787), .Y(register__n11650) );
  AO22x1_ASAP7_75t_R register___U3328 ( .A1(register__n9798), .A2(register__C6423_net61343), .B1(register__n10118), 
        .B2(register__net129787), .Y(register__n11420) );
  AO22x1_ASAP7_75t_R register___U3329 ( .A1(register__net91001), .A2(register__C6423_net61343), .B1(register__net89717), 
        .B2(register__net129787), .Y(register__n11289) );
  HB1xp67_ASAP7_75t_R register___U3330 ( .A(register__n11187), .Y(register__n4899) );
  AO22x1_ASAP7_75t_R register___U3331 ( .A1(register__n10495), .A2(register__net125426), .B1(register__n10450), .B2(
        net122862), .Y(register__n11187) );
  BUFx12f_ASAP7_75t_R register___U3332 ( .A(register__net140674), .Y(register__net64030) );
  BUFx6f_ASAP7_75t_R register___U3333 ( .A(register__net142400), .Y(register__net130838) );
  HB1xp67_ASAP7_75t_R register___U3334 ( .A(register__n12668), .Y(register__n4678) );
  NOR2xp67_ASAP7_75t_R register___U3335 ( .A(register__n2688), .B(register__n2687), .Y(register__n2686) );
  AND3x1_ASAP7_75t_R register___U3336 ( .A(register__n2947), .B(register__n7885), .C(register__n1076), .Y(register__n1043) );
  INVxp33_ASAP7_75t_R register___U3337 ( .A(register__n3710), .Y(register__n1815) );
  HB1xp67_ASAP7_75t_R register___U3338 ( .A(register__n13015), .Y(register__n4207) );
  BUFx6f_ASAP7_75t_R register___U3339 ( .A(register__net144162), .Y(register__net144689) );
  BUFx6f_ASAP7_75t_R register___U3340 ( .A(register__net143546), .Y(register__net144162) );
  HB1xp67_ASAP7_75t_R register___U3341 ( .A(register__n5604), .Y(register__n5603) );
  HB1xp67_ASAP7_75t_R register___U3342 ( .A(register__n12969), .Y(register__n2959) );
  INVx6_ASAP7_75t_R register___U3343 ( .A(register__n12071), .Y(register__n12058) );
  INVxp67_ASAP7_75t_R register___U3344 ( .A(register__n13166), .Y(register__n6403) );
  AND4x1_ASAP7_75t_R register___U3345 ( .A(register__n1511), .B(register__n12516), .C(register__n12511), .D(register__n12510), 
        .Y(register__n12512) );
  INVxp67_ASAP7_75t_R register___U3346 ( .A(register__n3891), .Y(register__n9404) );
  INVxp67_ASAP7_75t_R register___U3347 ( .A(register__n3432), .Y(register__n3997) );
  HB1xp67_ASAP7_75t_R register___U3348 ( .A(register__n3433), .Y(register__n3432) );
  OAI22xp33_ASAP7_75t_R register___U3349 ( .A1(register__n12111), .A2(register__n11863), .B1(register__n10305), .B2(
        n5341), .Y(register__n1015) );
  AND3x2_ASAP7_75t_R register___U3350 ( .A(register__n294), .B(WB_rd[2]), .C(register__n12488), .Y(
        n12485) );
  INVx2_ASAP7_75t_R register___U3351 ( .A(register__n12304), .Y(register__n12289) );
  INVx1_ASAP7_75t_R register___U3352 ( .A(register__n13290), .Y(register__n1016) );
  INVxp33_ASAP7_75t_R register___U3353 ( .A(register__n11873), .Y(register__n1819) );
  INVxp33_ASAP7_75t_R register___U3354 ( .A(register__n7633), .Y(register__n1807) );
  INVx1_ASAP7_75t_R register___U3355 ( .A(register__n12415), .Y(register__n12407) );
  INVx1_ASAP7_75t_R register___U3356 ( .A(register__n12852), .Y(register__n2271) );
  NOR2x1p5_ASAP7_75t_R register___U3357 ( .A(register__n2792), .B(register__n2791), .Y(register__n12852) );
  NOR2x2_ASAP7_75t_R register___U3358 ( .A(register__n12058), .B(register__n109), .Y(register__n2791) );
  INVx1_ASAP7_75t_R register___U3359 ( .A(register__n10975), .Y(register__n7675) );
  HB1xp67_ASAP7_75t_R register___U3360 ( .A(register__n12999), .Y(register__n4087) );
  HB1xp67_ASAP7_75t_R register___U3361 ( .A(register__n11699), .Y(register__n3117) );
  INVxp67_ASAP7_75t_R register___U3362 ( .A(register__n4411), .Y(register__n6740) );
  INVxp67_ASAP7_75t_R register___U3363 ( .A(register__n12607), .Y(register__n7255) );
  INVx1_ASAP7_75t_R register___U3364 ( .A(register__n13098), .Y(register__n1017) );
  INVx1_ASAP7_75t_R register___U3365 ( .A(register__n13311), .Y(register__n1018) );
  OAI22xp33_ASAP7_75t_R register___U3366 ( .A1(register__net63994), .A2(register__n11864), .B1(register__net89389), 
        .B2(register__n3680), .Y(register__n1020) );
  AOI22xp33_ASAP7_75t_R register___U3367 ( .A1(register__net64696), .A2(register__n1058), .B1(register__n7245), .B2(
        n1139), .Y(register__n13169) );
  INVx2_ASAP7_75t_R register___U3368 ( .A(register__net64704), .Y(register__net64672) );
  BUFx3_ASAP7_75t_R register___U3369 ( .A(register__n10640), .Y(register__n7245) );
  AOI22xp33_ASAP7_75t_R register___U3370 ( .A1(register__n12181), .A2(register__n1058), .B1(register__n1022), .B2(register__n103), 
        .Y(register__n13163) );
  CKINVDCx20_ASAP7_75t_R register___U3371 ( .A(register__n8728), .Y(register__n1022) );
  INVx2_ASAP7_75t_R register___U3372 ( .A(register__n12181), .Y(register__n12169) );
  BUFx4f_ASAP7_75t_R register___U3373 ( .A(register__net124704), .Y(register__net115027) );
  BUFx4f_ASAP7_75t_R register___U3374 ( .A(register__net99590), .Y(register__net117948) );
  HB1xp67_ASAP7_75t_R register___U3375 ( .A(register__n13017), .Y(register__n3433) );
  INVx1_ASAP7_75t_R register___U3376 ( .A(register__n13024), .Y(register__n1023) );
  CKINVDCx10_ASAP7_75t_R register___U3377 ( .A(n5), .Y(register__n12050) );
  BUFx3_ASAP7_75t_R register___U3378 ( .A(register__n10863), .Y(register__n4943) );
  AOI22xp33_ASAP7_75t_R register___U3379 ( .A1(register__n11987), .A2(register__n1058), .B1(register__n1024), .B2(register__n1140), .Y(register__n13174) );
  CKINVDCx20_ASAP7_75t_R register___U3380 ( .A(register__n9483), .Y(register__n1024) );
  INVx2_ASAP7_75t_R register___U3381 ( .A(register__n11987), .Y(register__n3666) );
  HB1xp67_ASAP7_75t_R register___U3382 ( .A(register__n8702), .Y(register__n4951) );
  NOR2xp67_ASAP7_75t_R register___U3383 ( .A(register__n969), .B(register__net89685), .Y(register__n5770) );
  CKINVDCx20_ASAP7_75t_R register___U3384 ( .A(register__n9481), .Y(register__n1026) );
  OAI22xp33_ASAP7_75t_R register___U3385 ( .A1(register__net64772), .A2(register__n187), .B1(register__net91001), .B2(
        n216), .Y(register__n1027) );
  INVx1_ASAP7_75t_R register___U3386 ( .A(register__n13256), .Y(register__n1028) );
  HB1xp67_ASAP7_75t_R register___U3387 ( .A(register__n5612), .Y(register__n5611) );
  INVxp67_ASAP7_75t_R register___U3388 ( .A(register__n13121), .Y(register__n4648) );
  BUFx12f_ASAP7_75t_R register___U3389 ( .A(register__n12245), .Y(register__n4966) );
  AND2x2_ASAP7_75t_R register___U3390 ( .A(register__n1770), .B(register__n11343), .Y(register__n1029) );
  AND2x2_ASAP7_75t_R register___U3391 ( .A(register__n11341), .B(register__n1029), .Y(register__n9175) );
  AND3x2_ASAP7_75t_R register___U3392 ( .A(register__n7597), .B(register__n1272), .C(register__n1769), .Y(register__n1030) );
  AND2x2_ASAP7_75t_R register___U3393 ( .A(register__n2828), .B(register__n1030), .Y(register__n11341) );
  BUFx12f_ASAP7_75t_R register___U3394 ( .A(register__n3690), .Y(register__n6465) );
  INVxp33_ASAP7_75t_R register___U3395 ( .A(register__n11814), .Y(register__n1777) );
  NOR2x1p5_ASAP7_75t_R register___U3396 ( .A(register__n1651), .B(register__n2707), .Y(register__n2709) );
  INVxp67_ASAP7_75t_R register___U3397 ( .A(register__n11812), .Y(register__n1632) );
  INVxp67_ASAP7_75t_R register___U3398 ( .A(register__n11300), .Y(register__n1031) );
  NOR2xp33_ASAP7_75t_R register___U3399 ( .A(register__net127626), .B(register__n11307), .Y(register__n1032) );
  NOR2xp33_ASAP7_75t_R register___U3400 ( .A(register__n1800), .B(register__n10642), .Y(register__n1034) );
  INVxp67_ASAP7_75t_R register___U3401 ( .A(register__n9513), .Y(register__n11307) );
  BUFx3_ASAP7_75t_R register___U3402 ( .A(register__C6422_net59756), .Y(register__net109872) );
  OAI22xp5_ASAP7_75t_R register___U3403 ( .A1(register__net66302), .A2(register__n8643), .B1(register__net64864), .B2(
        n1687), .Y(read_reg_data_2[5]) );
  HB1xp67_ASAP7_75t_R register___U3404 ( .A(register__C6423_net61326), .Y(register__n1035) );
  BUFx3_ASAP7_75t_R register___U3405 ( .A(register__C6423_net68950), .Y(register__net124706) );
  BUFx3_ASAP7_75t_R register___U3406 ( .A(register__C6423_net61326), .Y(register__net128121) );
  HB1xp67_ASAP7_75t_R register___U3407 ( .A(register__C6423_net68948), .Y(register__net136978) );
  HB1xp67_ASAP7_75t_R register___U3408 ( .A(register__net124706), .Y(register__net106379) );
  HB1xp67_ASAP7_75t_R register___U3409 ( .A(register__C6423_net68920), .Y(register__net106377) );
  HB1xp67_ASAP7_75t_R register___U3410 ( .A(register__net106377), .Y(register__C6423_net68930) );
  HB1xp67_ASAP7_75t_R register___U3411 ( .A(register__n11294), .Y(register__n5612) );
  OA22x2_ASAP7_75t_R register___U3412 ( .A1(register__net63322), .A2(register__n4033), .B1(register__n9734), .B2(register__n5050), 
        .Y(register__n12530) );
  NOR4xp75_ASAP7_75t_R register___U3413 ( .A(register__n1037), .B(register__n3236), .C(register__n2867), .D(register__n11471), 
        .Y(register__n11447) );
  CKINVDCx20_ASAP7_75t_R register___U3414 ( .A(register__n7259), .Y(register__n1037) );
  HB1xp67_ASAP7_75t_R register___U3415 ( .A(register__n11403), .Y(register__n4372) );
  OAI22xp5_ASAP7_75t_R register___U3416 ( .A1(register__net66308), .A2(register__n7021), .B1(register__n12164), .B2(
        n1687), .Y(read_reg_data_2[13]) );
  NOR2xp33_ASAP7_75t_R register___U3417 ( .A(register__n2565), .B(register__n2566), .Y(register__n2528) );
  INVx1_ASAP7_75t_R register___U3418 ( .A(register__n12711), .Y(register__n1038) );
  INVxp67_ASAP7_75t_R register___U3419 ( .A(register__net64802), .Y(register__net64768) );
  BUFx6f_ASAP7_75t_R register___U3420 ( .A(register__net147378), .Y(register__C6423_net74857) );
  INVxp67_ASAP7_75t_R register___U3421 ( .A(register__n2117), .Y(register__n1659) );
  INVxp33_ASAP7_75t_R register___U3422 ( .A(register__n1657), .Y(register__n1661) );
  INVxp33_ASAP7_75t_R register___U3423 ( .A(register__n2117), .Y(register__n1660) );
  INVx2_ASAP7_75t_R register___U3424 ( .A(register__n2121), .Y(register__n2122) );
  HB1xp67_ASAP7_75t_R register___U3425 ( .A(register__n3961), .Y(register__n3960) );
  INVx2_ASAP7_75t_R register___U3426 ( .A(register__n1136), .Y(register__n1141) );
  NOR3xp33_ASAP7_75t_R register___U3427 ( .A(register__n9231), .B(register__n1041), .C(register__n1042), .Y(register__n1040) );
  OAI22xp33_ASAP7_75t_R register___U3428 ( .A1(register__n420), .A2(register__n7098), .B1(register__n801), .B2(register__n8589), 
        .Y(register__n1042) );
  INVx1_ASAP7_75t_R register___U3429 ( .A(register__n1947), .Y(register__n1948) );
  INVx1_ASAP7_75t_R register___U3430 ( .A(register__n2105), .Y(register__n2106) );
  INVxp67_ASAP7_75t_R register___U3431 ( .A(register__n12658), .Y(register__n7076) );
  AND2x2_ASAP7_75t_R register___U3432 ( .A(register__n3118), .B(register__n1043), .Y(register__n11678) );
  INVx1_ASAP7_75t_R register___U3433 ( .A(register__n11698), .Y(register__n2947) );
  BUFx2_ASAP7_75t_R register___U3434 ( .A(register__n7886), .Y(register__n3118) );
  INVx6_ASAP7_75t_R register___U3435 ( .A(register__n3378), .Y(register__n12115) );
  BUFx12f_ASAP7_75t_R register___U3436 ( .A(register__n3366), .Y(register__n3378) );
  INVx1_ASAP7_75t_R register___U3437 ( .A(register__n13331), .Y(register__n1044) );
  HB1xp67_ASAP7_75t_R register___U3438 ( .A(register__n1382), .Y(register__net145264) );
  INVx3_ASAP7_75t_R register___U3439 ( .A(register__net64964), .Y(register__net64920) );
  INVxp67_ASAP7_75t_R register___U3440 ( .A(register__n5763), .Y(register__n7902) );
  BUFx2_ASAP7_75t_R register___U3441 ( .A(register__n3237), .Y(register__n3236) );
  CKINVDCx12_ASAP7_75t_R register___U3442 ( .A(n7), .Y(register__net128430) );
  OAI22xp5_ASAP7_75t_R register___U3443 ( .A1(register__net66314), .A2(register__n7614), .B1(register__net126178), .B2(
        n1687), .Y(read_reg_data_2[23]) );
  INVxp67_ASAP7_75t_R register___U3444 ( .A(register__n4427), .Y(register__n5217) );
  OAI22xp33_ASAP7_75t_R register___U3445 ( .A1(register__n12196), .A2(register__n1137), .B1(register__n8718), .B2(register__n1147), .Y(register__n1748) );
  HB1xp67_ASAP7_75t_R register___U3446 ( .A(register__n4412), .Y(register__n4411) );
  AO22x1_ASAP7_75t_R register___U3447 ( .A1(register__n9816), .A2(register__net93569), .B1(register__n10227), .B2(
        net147378), .Y(register__n11384) );
  AO22x1_ASAP7_75t_R register___U3448 ( .A1(register__n8347), .A2(register__net93569), .B1(register__n8803), .B2(
        net147378), .Y(register__n11470) );
  AO22x1_ASAP7_75t_R register___U3449 ( .A1(register__n5645), .A2(register__n1106), .B1(register__n6039), .B2(register__n285), 
        .Y(register__n11217) );
  AO22x1_ASAP7_75t_R register___U3450 ( .A1(register__net116361), .A2(register__net93569), .B1(register__net112729), 
        .B2(register__n284), .Y(register__n11295) );
  OAI22xp5_ASAP7_75t_R register___U3451 ( .A1(register__n54), .A2(register__n7323), .B1(register__net61369), .B2(register__n12033), .Y(read_reg_data_1[3]) );
  AND3x1_ASAP7_75t_R register___U3452 ( .A(register__n1582), .B(register__n7596), .C(register__n3792), .Y(register__n7593) );
  INVx2_ASAP7_75t_R register___U3453 ( .A(register__n11228), .Y(register__n7063) );
  NAND3x1_ASAP7_75t_R register___U3454 ( .A(register__n8225), .B(register__n269), .C(register__n5916), .Y(register__n1048) );
  BUFx6f_ASAP7_75t_R register___U3455 ( .A(register__net141041), .Y(register__net143489) );
  BUFx6f_ASAP7_75t_R register___U3456 ( .A(register__net91921), .Y(register__net141041) );
  NOR2xp33_ASAP7_75t_R register___U3457 ( .A(register__net89209), .B(register__n1161), .Y(register__n6397) );
  XNOR2xp5_ASAP7_75t_R register___U3458 ( .A(register__n244), .B(register__n717), .Y(register__n12511) );
  BUFx3_ASAP7_75t_R register___U3459 ( .A(register__n3339), .Y(register__n3296) );
  HB1xp67_ASAP7_75t_R register___U3460 ( .A(register__n2886), .Y(register__n2856) );
  BUFx3_ASAP7_75t_R register___U3461 ( .A(register__n3296), .Y(register__n2835) );
  BUFx6f_ASAP7_75t_R register___U3462 ( .A(register__n3295), .Y(register__n11744) );
  INVx3_ASAP7_75t_R register___U3463 ( .A(register__n3339), .Y(register__n3337) );
  INVxp67_ASAP7_75t_R register___U3464 ( .A(register__n5000), .Y(register__n7074) );
  HB1xp67_ASAP7_75t_R register___U3465 ( .A(register__n5001), .Y(register__n5000) );
  HB1xp67_ASAP7_75t_R register___U3466 ( .A(register__n12655), .Y(register__n5001) );
  AO22x1_ASAP7_75t_R register___U3467 ( .A1(register__n7705), .A2(register__n85), .B1(register__n8031), .B2(register__n422), .Y(
        n11574) );
  AO22x1_ASAP7_75t_R register___U3468 ( .A1(register__n9710), .A2(register__n85), .B1(register__n10040), .B2(
        C6423_net61335), .Y(register__n11442) );
  AO22x1_ASAP7_75t_R register___U3469 ( .A1(register__n7539), .A2(register__n85), .B1(register__n10323), .B2(register__n2086), 
        .Y(register__n11652) );
  AO22x1_ASAP7_75t_R register___U3470 ( .A1(register__n9832), .A2(register__n85), .B1(register__n10128), .B2(register__n422), .Y(
        n11594) );
  AO22x1_ASAP7_75t_R register___U3471 ( .A1(register__net90729), .A2(register__n85), .B1(register__net89813), .B2(register__n422), 
        .Y(register__n11272) );
  AO22x1_ASAP7_75t_R register___U3472 ( .A1(register__n9700), .A2(register__n85), .B1(register__n10050), .B2(
        C6423_net61335), .Y(register__n11168) );
  AO22x1_ASAP7_75t_R register___U3473 ( .A1(register__n9053), .A2(register__n85), .B1(register__n8375), .B2(
        C6423_net61335), .Y(register__n11694) );
  AND2x2_ASAP7_75t_R register___U3474 ( .A(rs2[1]), .B(rs2[0]), 
        .Y(register__n7052) );
  HB1xp67_ASAP7_75t_R register___U3475 ( .A(register__n12141), .Y(register__n4635) );
  BUFx2_ASAP7_75t_R register___U3476 ( .A(register__n3543), .Y(register__n3917) );
  INVx1_ASAP7_75t_R register___U3477 ( .A(register__n3299), .Y(register__n12374) );
  INVx2_ASAP7_75t_R register___U3478 ( .A(register__n12374), .Y(register__n1880) );
  BUFx12f_ASAP7_75t_R register___U3479 ( .A(register__n12416), .Y(register__n3726) );
  HB1xp67_ASAP7_75t_R register___U3480 ( .A(register__n3726), .Y(register__n12415) );
  INVx1_ASAP7_75t_R register___U3481 ( .A(register__n12696), .Y(register__n1051) );
  CKINVDCx20_ASAP7_75t_R register___U3482 ( .A(register__n9597), .Y(register__n1052) );
  HB1xp67_ASAP7_75t_R register___U3483 ( .A(register__n11469), .Y(register__n3237) );
  AO22x1_ASAP7_75t_R register___U3484 ( .A1(register__n9855), .A2(register__n1105), .B1(register__n10281), .B2(register__n285), 
        .Y(register__n11636) );
  INVxp67_ASAP7_75t_R register___U3485 ( .A(register__n13258), .Y(register__n7287) );
  HB1xp67_ASAP7_75t_R register___U3486 ( .A(register__n4428), .Y(register__n4427) );
  NOR2xp67_ASAP7_75t_R register___U3487 ( .A(register__n12061), .B(register__n4035), .Y(register__n2793) );
  AOI22xp33_ASAP7_75t_R register___U3488 ( .A1(register__net62708), .A2(register__n1586), .B1(register__n1053), .B2(
        n2935), .Y(register__n12691) );
  CKINVDCx20_ASAP7_75t_R register___U3489 ( .A(register__n7847), .Y(register__n1053) );
  INVx2_ASAP7_75t_R register___U3490 ( .A(register__n3022), .Y(register__n1586) );
  INVx1_ASAP7_75t_R register___U3491 ( .A(register__n13059), .Y(register__n1054) );
  INVxp67_ASAP7_75t_R register___U3492 ( .A(register__net64804), .Y(register__net64770) );
  BUFx6f_ASAP7_75t_R register___U3493 ( .A(register__net64802), .Y(register__net138526) );
  HB1xp67_ASAP7_75t_R register___U3494 ( .A(register__n5764), .Y(register__n5763) );
  AO22x1_ASAP7_75t_R register___U3495 ( .A1(register__n9642), .A2(register__net109849), .B1(register__n9969), .B2(register__n645), 
        .Y(register__n11579) );
  AO22x1_ASAP7_75t_R register___U3496 ( .A1(register__n9650), .A2(register__n481), .B1(register__n9977), .B2(register__n648), .Y(
        n11259) );
  AO22x1_ASAP7_75t_R register___U3497 ( .A1(register__n10440), .A2(register__n481), .B1(register__n10469), .B2(register__n539), 
        .Y(register__n11516) );
  AO22x1_ASAP7_75t_R register___U3498 ( .A1(register__n9656), .A2(register__n481), .B1(register__n9983), .B2(register__n638), .Y(
        n11194) );
  AO22x1_ASAP7_75t_R register___U3499 ( .A1(register__n9887), .A2(register__n481), .B1(register__n10311), .B2(
        C6423_net61348), .Y(register__n11471) );
  AO22x1_ASAP7_75t_R register___U3500 ( .A1(register__n8807), .A2(register__n482), .B1(register__n8817), .B2(
        C6423_net61348), .Y(register__n11559) );
  AO22x1_ASAP7_75t_R register___U3501 ( .A1(register__n8127), .A2(register__n482), .B1(register__n10467), .B2(
        C6423_net61348), .Y(register__n11725) );
  AO22x1_ASAP7_75t_R register___U3502 ( .A1(register__n9672), .A2(register__n1950), .B1(register__n9919), .B2(register__n767), 
        .Y(register__n11535) );
  AO22x1_ASAP7_75t_R register___U3503 ( .A1(register__n9726), .A2(register__n2004), .B1(register__n5679), .B2(register__n767), 
        .Y(register__n11315) );
  AO22x1_ASAP7_75t_R register___U3504 ( .A1(register__n1967), .A2(register__n6974), .B1(register__n10473), .B2(register__n767), 
        .Y(register__n11653) );
  AO22x1_ASAP7_75t_R register___U3505 ( .A1(register__n9678), .A2(register__n1967), .B1(register__n9925), .B2(register__n767), 
        .Y(register__n11214) );
  AO22x1_ASAP7_75t_R register___U3506 ( .A1(register__n10436), .A2(register__n1966), .B1(register__n10475), .B2(register__n767), 
        .Y(register__n11673) );
  AO22x1_ASAP7_75t_R register___U3507 ( .A1(register__n9758), .A2(register__n1967), .B1(register__n8491), .B2(register__n767), 
        .Y(register__n11423) );
  AO22x1_ASAP7_75t_R register___U3508 ( .A1(register__net90833), .A2(register__n1967), .B1(register__net90149), .B2(
        n767), .Y(register__n11292) );
  AO22x1_ASAP7_75t_R register___U3509 ( .A1(register__n9337), .A2(register__n1967), .B1(register__n8783), .B2(register__n767), 
        .Y(register__n11336) );
  AO22x1_ASAP7_75t_R register___U3510 ( .A1(register__n7573), .A2(register__n1967), .B1(register__n10297), .B2(register__n767), 
        .Y(register__n11718) );
  HB1xp67_ASAP7_75t_R register___U3511 ( .A(register__n11695), .Y(register__n5604) );
  AO22x1_ASAP7_75t_R register___U3512 ( .A1(register__net90545), .A2(register__n1967), .B1(register__net89037), .B2(
        n767), .Y(register__n11612) );
  AO22x1_ASAP7_75t_R register___U3513 ( .A1(register__n9756), .A2(register__C6423_net61333), .B1(register__n9062), .B2(
        C6423_net61331), .Y(register__n11695) );
  INVx1_ASAP7_75t_R register___U3514 ( .A(register__n13330), .Y(register__n1055) );
  BUFx12f_ASAP7_75t_R register___U3515 ( .A(register__net73061), .Y(register__net104559) );
  BUFx12f_ASAP7_75t_R register___U3516 ( .A(register__n3570), .Y(register__n3532) );
  AO22x1_ASAP7_75t_R register___U3517 ( .A1(register__n5443), .A2(register__n3336), .B1(register__n1754), .B2(register__n1266), 
        .Y(register__n1753) );
  INVxp33_ASAP7_75t_R register___U3518 ( .A(register__n1753), .Y(register__n13131) );
  AO22x1_ASAP7_75t_R register___U3519 ( .A1(register__n12183), .A2(register__n88), .B1(register__n1057), .B2(register__n1713), 
        .Y(register__n1056) );
  CKINVDCx20_ASAP7_75t_R register___U3520 ( .A(register__n10205), .Y(register__n1057) );
  HB1xp67_ASAP7_75t_R register___U3521 ( .A(register__n12638), .Y(register__n4412) );
  HB1xp67_ASAP7_75t_R register___U3522 ( .A(register__n13156), .Y(register__n3739) );
  AO22x1_ASAP7_75t_R register___U3523 ( .A1(register__n8813), .A2(register__net129747), .B1(register__n8821), .B2(
        net123857), .Y(register__n11048) );
  AO22x1_ASAP7_75t_R register___U3524 ( .A1(register__n9686), .A2(register__C6422_net60422), .B1(register__n9957), .B2(
        net123857), .Y(register__n10922) );
  BUFx12f_ASAP7_75t_R register___U3525 ( .A(register__n3600), .Y(register__n3599) );
  BUFx12f_ASAP7_75t_R register___U3526 ( .A(register__n3381), .Y(register__n5499) );
  HB1xp67_ASAP7_75t_R register___U3527 ( .A(register__n13169), .Y(register__n3827) );
  HB1xp67_ASAP7_75t_R register___U3528 ( .A(register__n13173), .Y(register__n3741) );
  HB1xp67_ASAP7_75t_R register___U3529 ( .A(register__n13174), .Y(register__n3825) );
  HB1xp67_ASAP7_75t_R register___U3530 ( .A(register__n13161), .Y(register__n3961) );
  HB1xp67_ASAP7_75t_R register___U3531 ( .A(register__n13163), .Y(register__n3969) );
  AO21x1_ASAP7_75t_R register___U3532 ( .A1(register__net91375), .A2(register__net114704), .B(register__n1059), .Y(
        n2619) );
  AND2x2_ASAP7_75t_R register___U3533 ( .A(register__n1116), .B(register__n2633), .Y(register__n1059) );
  AO22x1_ASAP7_75t_R register___U3534 ( .A1(register__n9901), .A2(register__n309), .B1(register__n10333), .B2(register__n284), 
        .Y(register__n11676) );
  AO22x1_ASAP7_75t_R register___U3535 ( .A1(register__net91069), .A2(register__net93569), .B1(register__net89909), .B2(
        n284), .Y(register__n11276) );
  INVxp33_ASAP7_75t_R register___U3536 ( .A(register__n4851), .Y(register__n1847) );
  INVxp33_ASAP7_75t_R register___U3537 ( .A(register__n4851), .Y(register__n1844) );
  INVxp33_ASAP7_75t_R register___U3538 ( .A(register__n4851), .Y(register__n1846) );
  INVxp33_ASAP7_75t_R register___U3539 ( .A(register__n4851), .Y(register__n1845) );
  AO22x1_ASAP7_75t_R register___U3540 ( .A1(register__n6669), .A2(register__n920), .B1(register__n10315), .B2(register__net150890), .Y(register__n11469) );
  AOI22xp33_ASAP7_75t_R register___U3541 ( .A1(register__n12066), .A2(register__n1146), .B1(register__n1060), .B2(register__n103), 
        .Y(register__n13168) );
  CKINVDCx20_ASAP7_75t_R register___U3542 ( .A(register__n8720), .Y(register__n1060) );
  AOI22xp33_ASAP7_75t_R register___U3543 ( .A1(register__n9409), .A2(register__net122599), .B1(register__n9423), .B2(
        C6423_net68766), .Y(register__n1061) );
  INVxp67_ASAP7_75t_R register___U3544 ( .A(register__n12581), .Y(register__n7904) );
  INVx2_ASAP7_75t_R register___U3545 ( .A(register__n1971), .Y(register__n1540) );
  INVx2_ASAP7_75t_R register___U3546 ( .A(register__n5957), .Y(register__n6830) );
  AO22x1_ASAP7_75t_R register___U3547 ( .A1(register__net88412), .A2(register__n413), .B1(register__net88628), .B2(
        net126602), .Y(register__n10807) );
  AO22x1_ASAP7_75t_R register___U3548 ( .A1(register__n8763), .A2(register__n413), .B1(register__n9359), .B2(
        C6422_net60401), .Y(register__n10558) );
  NAND2xp33_ASAP7_75t_R register___U3549 ( .A(register__net131638), .B(register__n2524), .Y(register__n2511) );
  NAND2xp33_ASAP7_75t_R register___U3550 ( .A(register__net131638), .B(register__net106200), .Y(register__n2616) );
  HB1xp67_ASAP7_75t_R register___U3551 ( .A(register__n12637), .Y(register__n4428) );
  INVxp33_ASAP7_75t_R register___U3552 ( .A(register__net130482), .Y(register__n1657) );
  OAI22xp33_ASAP7_75t_R register___U3553 ( .A1(register__n12429), .A2(register__n2826), .B1(register__n10383), .B2(
        n1933), .Y(register__n1062) );
  BUFx2_ASAP7_75t_R register___U3554 ( .A(register__n11925), .Y(register__n3373) );
  INVxp67_ASAP7_75t_R register___U3555 ( .A(register__n11938), .Y(register__n11925) );
  AOI22xp33_ASAP7_75t_R register___U3556 ( .A1(register__n12442), .A2(register__n11783), .B1(register__n1063), .B2(
        n1576), .Y(register__n12891) );
  CKINVDCx20_ASAP7_75t_R register___U3557 ( .A(register__n10425), .Y(register__n1063) );
  INVx1_ASAP7_75t_R register___U3558 ( .A(register__n12834), .Y(register__n1064) );
  INVx1_ASAP7_75t_R register___U3559 ( .A(register__n12803), .Y(register__n1065) );
  NOR2xp33_ASAP7_75t_R register___U3560 ( .A(register__n1420), .B(register__n1066), .Y(register__n1067) );
  NOR2xp33_ASAP7_75t_R register___U3561 ( .A(register__n1067), .B(register__n2682), .Y(register__n2683) );
  INVxp33_ASAP7_75t_R register___U3562 ( .A(register__net89041), .Y(register__n1066) );
  BUFx3_ASAP7_75t_R register___U3563 ( .A(register__net107870), .Y(register__net89041) );
  NOR4xp25_ASAP7_75t_R register___U3564 ( .A(register__n1230), .B(register__n10540), .C(register__n10541), .D(register__n10542), 
        .Y(register__n10523) );
  INVx1_ASAP7_75t_R register___U3565 ( .A(register__n6416), .Y(register__n1230) );
  HB1xp67_ASAP7_75t_R register___U3566 ( .A(register__n12494), .Y(register__n4579) );
  HB1xp67_ASAP7_75t_R register___U3567 ( .A(register__n11485), .Y(register__n5626) );
  AO22x1_ASAP7_75t_R register___U3568 ( .A1(register__n9384), .A2(register__n883), .B1(register__n9380), .B2(register__net122862), 
        .Y(register__n11485) );
  INVx6_ASAP7_75t_R register___U3569 ( .A(register__n12389), .Y(register__n12377) );
  INVx1_ASAP7_75t_R register___U3570 ( .A(register__n10550), .Y(register__n7670) );
  INVxp67_ASAP7_75t_R register___U3571 ( .A(register__n5968), .Y(register__n8238) );
  AOI22xp33_ASAP7_75t_R register___U3572 ( .A1(register__n12387), .A2(register__n82), .B1(register__n1068), .B2(register__n2801), 
        .Y(register__n12809) );
  AO21x2_ASAP7_75t_R register___U3573 ( .A1(register__net90665), .A2(register__net125426), .B(register__n2618), .Y(
        n1070) );
  NOR2x1_ASAP7_75t_R register___U3574 ( .A(register__n1070), .B(register__n2619), .Y(register__n2620) );
  BUFx6f_ASAP7_75t_R register___U3575 ( .A(register__net112407), .Y(register__net90665) );
  OAI21xp33_ASAP7_75t_R register___U3576 ( .A1(register__C6423_net60775), .A2(register__n714), .B(register__n2617), .Y(
        n2618) );
  INVxp67_ASAP7_75t_R register___U3577 ( .A(register__n11288), .Y(register__n1071) );
  AO22x1_ASAP7_75t_R register___U3578 ( .A1(register__n9867), .A2(register__C6422_net60415), .B1(register__n10291), 
        .B2(register__net88727), .Y(register__n11029) );
  AO22x1_ASAP7_75t_R register___U3579 ( .A1(register__net93797), .A2(register__C6422_net60415), .B1(register__net115999), .B2(register__net88727), .Y(register__n10813) );
  OAI22x1_ASAP7_75t_R register___U3580 ( .A1(register__net63320), .A2(register__n1989), .B1(register__n10268), .B2(
        n11852), .Y(register__n1072) );
  INVx4_ASAP7_75t_R register___U3581 ( .A(register__n4728), .Y(register__n12395) );
  INVxp67_ASAP7_75t_R register___U3582 ( .A(register__n3688), .Y(register__n7632) );
  HB1xp67_ASAP7_75t_R register___U3583 ( .A(register__n3689), .Y(register__n3688) );
  OAI21xp33_ASAP7_75t_R register___U3584 ( .A1(register__n2585), .A2(register__net66306), .B(register__n2589), .Y(
        read_reg_data_2[11]) );
  BUFx6f_ASAP7_75t_R register___U3585 ( .A(register__net117889), .Y(register__net125797) );
  HB1xp67_ASAP7_75t_R register___U3586 ( .A(register__net125797), .Y(register__net128105) );
  HB1xp67_ASAP7_75t_R register___U3587 ( .A(register__net128105), .Y(register__C6423_net69560) );
  AOI22xp33_ASAP7_75t_R register___U3588 ( .A1(register__net147378), .A2(register__net88548), .B1(register__net93569), 
        .B2(register__net88472), .Y(register__n2456) );
  INVx1_ASAP7_75t_R register___U3589 ( .A(register__n12756), .Y(register__n1075) );
  BUFx3_ASAP7_75t_R register___U3590 ( .A(register__n12450), .Y(register__n6267) );
  INVx1_ASAP7_75t_R register___U3591 ( .A(register__n11697), .Y(register__n1076) );
  INVx1_ASAP7_75t_R register___U3592 ( .A(register__n12726), .Y(register__n1077) );
  INVx1_ASAP7_75t_R register___U3593 ( .A(register__n13276), .Y(register__n1078) );
  BUFx12f_ASAP7_75t_R register___U3594 ( .A(register__n3341), .Y(register__n12389) );
  INVxp67_ASAP7_75t_R register___U3595 ( .A(register__n3609), .Y(register__n5547) );
  INVxp67_ASAP7_75t_R register___U3596 ( .A(register__n4208), .Y(register__n7286) );
  HB1xp67_ASAP7_75t_R register___U3597 ( .A(register__n4209), .Y(register__n4208) );
  AO22x1_ASAP7_75t_R register___U3598 ( .A1(register__n3536), .A2(register__n5721), .B1(register__n1410), .B2(register__n1411), 
        .Y(register__n1079) );
  BUFx6f_ASAP7_75t_R register___U3599 ( .A(register__n3512), .Y(register__n5041) );
  AO22x1_ASAP7_75t_R register___U3600 ( .A1(register__net90965), .A2(register__net110414), .B1(register__net89689), 
        .B2(register__n1074), .Y(register__n11293) );
  HB1xp67_ASAP7_75t_R register___U3601 ( .A(register__net100798), .Y(register__net62694) );
  INVxp67_ASAP7_75t_R register___U3602 ( .A(register__n12586), .Y(register__n4383) );
  HB1xp67_ASAP7_75t_R register___U3603 ( .A(register__n11468), .Y(register__n3235) );
  AO22x1_ASAP7_75t_R register___U3604 ( .A1(register__n9750), .A2(register__net110414), .B1(register__n10126), .B2(
        n1074), .Y(register__n11402) );
  BUFx12f_ASAP7_75t_R register___U3605 ( .A(register__net125327), .Y(register__net129617) );
  HB1xp67_ASAP7_75t_R register___U3606 ( .A(register__n3181), .Y(register__n3180) );
  BUFx3_ASAP7_75t_R register___U3607 ( .A(register__n12355), .Y(register__n3346) );
  INVx2_ASAP7_75t_R register___U3608 ( .A(register__net62708), .Y(register__net62672) );
  BUFx3_ASAP7_75t_R register___U3609 ( .A(register__net141985), .Y(register__net62708) );
  BUFx6f_ASAP7_75t_R register___U3610 ( .A(register__n6267), .Y(register__n12441) );
  HB1xp67_ASAP7_75t_R register___U3611 ( .A(register__n5232), .Y(register__n4119) );
  INVxp33_ASAP7_75t_R register___U3612 ( .A(register__n4117), .Y(register__n5232) );
  BUFx6f_ASAP7_75t_R register___U3613 ( .A(register__net73055), .Y(register__net129518) );
  INVx2_ASAP7_75t_R register___U3614 ( .A(register__net129518), .Y(register__n1680) );
  BUFx3_ASAP7_75t_R register___U3615 ( .A(register__net129518), .Y(register__net127289) );
  INVx1_ASAP7_75t_R register___U3616 ( .A(register__net129518), .Y(register__n2111) );
  INVxp67_ASAP7_75t_R register___U3617 ( .A(register__n12831), .Y(register__n8595) );
  INVxp67_ASAP7_75t_R register___U3618 ( .A(register__n6252), .Y(register__n6996) );
  AO22x1_ASAP7_75t_R register___U3619 ( .A1(register__n8755), .A2(register__C6423_net61326), .B1(register__n10060), 
        .B2(register__n1999), .Y(register__n11228) );
  NOR2xp33_ASAP7_75t_R register___U3620 ( .A(register__C6423_net60882), .B(register__n1995), .Y(register__n2691) );
  CKINVDCx10_ASAP7_75t_R register___U3621 ( .A(write_data[28]), .Y(register__n12450) );
  NOR3x1_ASAP7_75t_R register___U3622 ( .A(register__n1082), .B(register__n2274), .C(register__n5336), .Y(register__n7941) );
  HB1xp67_ASAP7_75t_R register___U3623 ( .A(register__net131654), .Y(register__n1964) );
  INVx2_ASAP7_75t_R register___U3624 ( .A(register__n12525), .Y(register__n6689) );
  INVx6_ASAP7_75t_R register___U3625 ( .A(register__n12446), .Y(register__n12430) );
  BUFx6f_ASAP7_75t_R register___U3626 ( .A(register__n4634), .Y(register__n12130) );
  INVxp33_ASAP7_75t_R register___U3627 ( .A(register__n11669), .Y(register__n1084) );
  HB1xp67_ASAP7_75t_R register___U3628 ( .A(register__n4278), .Y(register__n4156) );
  BUFx6f_ASAP7_75t_R register___U3629 ( .A(register__n7258), .Y(register__n3454) );
  INVx2_ASAP7_75t_R register___U3630 ( .A(register__n3481), .Y(register__n12434) );
  BUFx6f_ASAP7_75t_R register___U3631 ( .A(register__n3454), .Y(register__n3481) );
  INVx2_ASAP7_75t_R register___U3632 ( .A(register__net64872), .Y(register__net64840) );
  BUFx2_ASAP7_75t_R register___U3633 ( .A(register__net143364), .Y(register__net64872) );
  HB1xp67_ASAP7_75t_R register___U3634 ( .A(register__n5182), .Y(register__n3390) );
  INVx3_ASAP7_75t_R register___U3635 ( .A(register__n12410), .Y(register__n12396) );
  INVx1_ASAP7_75t_R register___U3636 ( .A(register__n12746), .Y(register__n1086) );
  AND2x2_ASAP7_75t_R register___U3637 ( .A(register__n1087), .B(register__n1088), .Y(register__n12746) );
  AND3x2_ASAP7_75t_R register___U3638 ( .A(register__n5247), .B(WB_rd[3]), .C(RegWrite), 
        .Y(register__n12495) );
  INVxp33_ASAP7_75t_R register___U3639 ( .A(register__n10297), .Y(register__n1238) );
  INVx1_ASAP7_75t_R register___U3640 ( .A(register__n12749), .Y(register__n8625) );
  INVx4_ASAP7_75t_R register___U3641 ( .A(register__n3482), .Y(register__n12431) );
  BUFx12f_ASAP7_75t_R register___U3642 ( .A(register__n3455), .Y(register__n3482) );
  INVx3_ASAP7_75t_R register___U3643 ( .A(register__n12133), .Y(register__n12112) );
  INVxp33_ASAP7_75t_R register___U3644 ( .A(register__n3569), .Y(register__n2234) );
  BUFx12_ASAP7_75t_R register___U3645 ( .A(register__net145523), .Y(register__net145772) );
  OAI22xp5_ASAP7_75t_R register___U3646 ( .A1(register__n53), .A2(register__n9179), .B1(register__net61369), .B2(register__n12133), .Y(read_reg_data_1[12]) );
  INVxp67_ASAP7_75t_R register___U3647 ( .A(register__n6025), .Y(register__n9208) );
  HB1xp67_ASAP7_75t_R register___U3648 ( .A(register__n6026), .Y(register__n6025) );
  NAND2x1_ASAP7_75t_R register___U3649 ( .A(register__n4913), .B(register__n2798), .Y(register__n2262) );
  AO22x1_ASAP7_75t_R register___U3650 ( .A1(register__n9301), .A2(register__n77), .B1(register__n10337), .B2(register__n75), .Y(
        n11075) );
  NAND2x1p5_ASAP7_75t_R register___U3651 ( .A(register__n2516), .B(register__n2518), .Y(register__n2517) );
  AND2x2_ASAP7_75t_R register___U3652 ( .A(register__register__n6999), .B(register__n6), .Y(register__n1089) );
  AND3x1_ASAP7_75t_R register___U3653 ( .A(register__n1089), .B(register__n9152), .C(register__n6998), .Y(register__n10655) );
  INVx1_ASAP7_75t_R register___U3654 ( .A(register__n5274), .Y(register__n6998) );
  INVxp67_ASAP7_75t_R register___U3655 ( .A(register__n4497), .Y(register__n6173) );
  HB1xp67_ASAP7_75t_R register___U3656 ( .A(register__n4498), .Y(register__n4497) );
  HB1xp67_ASAP7_75t_R register___U3657 ( .A(register__n12364), .Y(register__n3265) );
  HB1xp67_ASAP7_75t_R register___U3658 ( .A(register__n11368), .Y(register__n6026) );
  INVxp67_ASAP7_75t_R register___U3659 ( .A(register__n1949), .Y(register__n1551) );
  BUFx6f_ASAP7_75t_R register___U3660 ( .A(register__net63222), .Y(register__net143546) );
  HB1xp67_ASAP7_75t_R register___U3661 ( .A(register__n3456), .Y(register__n4036) );
  INVx1_ASAP7_75t_R register___U3662 ( .A(register__n13076), .Y(register__n1091) );
  XNOR2xp5_ASAP7_75t_R register___U3663 ( .A(register__n1011), .B(register__n4264), .Y(register__n12510) );
  BUFx12f_ASAP7_75t_R register___U3664 ( .A(register__n3670), .Y(register__n3669) );
  BUFx6f_ASAP7_75t_R register___U3665 ( .A(register__n3455), .Y(register__n12444) );
  HB1xp67_ASAP7_75t_R register___U3666 ( .A(register__n13180), .Y(register__n4410) );
  NAND2xp5_ASAP7_75t_R register___U3667 ( .A(register__n9353), .B(register__n1226), .Y(register__n1093) );
  NAND2xp33_ASAP7_75t_R register___U3668 ( .A(register__n8793), .B(register__n75), .Y(register__n1094) );
  NAND2xp33_ASAP7_75t_R register___U3669 ( .A(register__n1093), .B(register__n1094), .Y(register__n11052) );
  HB1xp67_ASAP7_75t_R register___U3670 ( .A(register__n11052), .Y(register__n5606) );
  BUFx3_ASAP7_75t_R register___U3671 ( .A(register__n12425), .Y(register__n3304) );
  OAI22xp5_ASAP7_75t_R register___U3672 ( .A1(register__n54), .A2(register__n7273), .B1(register__net61369), .B2(register__n12178), .Y(read_reg_data_1[14]) );
  OAI22xp33_ASAP7_75t_R register___U3673 ( .A1(register__n11922), .A2(register__n337), .B1(register__n9634), .B2(register__n345), 
        .Y(register__n1096) );
  CKINVDCx20_ASAP7_75t_R register___U3674 ( .A(register__net90109), .Y(register__n1097) );
  OAI22xp33_ASAP7_75t_R register___U3675 ( .A1(register__n11922), .A2(register__n699), .B1(register__n9501), .B2(register__n678), 
        .Y(register__n1099) );
  INVx6_ASAP7_75t_R register___U3676 ( .A(register__net145522), .Y(register__net64850) );
  AO22x1_ASAP7_75t_R register___U3677 ( .A1(register__net64964), .A2(register__n5531), .B1(register__n1102), .B2(register__n1120), 
        .Y(register__n1101) );
  CKINVDCx20_ASAP7_75t_R register___U3678 ( .A(register__n9260), .Y(register__n1102) );
  OAI22x1_ASAP7_75t_R register___U3679 ( .A1(register__net64916), .A2(register__n1989), .B1(register__n8082), .B2(register__n2961), .Y(register__n1103) );
  HB1xp67_ASAP7_75t_R register___U3680 ( .A(register__n5182), .Y(register__n3170) );
  NOR2xp33_ASAP7_75t_R register___U3681 ( .A(register__n2013), .B(register__n2690), .Y(register__n2692) );
  HB1xp67_ASAP7_75t_R register___U3682 ( .A(register__n12633), .Y(register__n5764) );
  INVxp67_ASAP7_75t_R register___U3683 ( .A(register__n3430), .Y(register__n5236) );
  NAND3xp33_ASAP7_75t_R register___U3684 ( .A(register__n564), .B(register__n849), .C(register__n1422), .Y(register__n1104) );
  BUFx6f_ASAP7_75t_R register___U3685 ( .A(register__n12130), .Y(register__n3379) );
  HB1xp67_ASAP7_75t_R register___U3686 ( .A(register__n12770), .Y(register__n4498) );
  NOR2xp33_ASAP7_75t_R register___U3687 ( .A(register__n1335), .B(register__n7697), .Y(register__n1105) );
  HB1xp67_ASAP7_75t_R register___U3688 ( .A(register__n309), .Y(register__C6423_net74825) );
  HB1xp67_ASAP7_75t_R register___U3689 ( .A(register__C6423_net74825), .Y(register__net146317) );
  INVxp67_ASAP7_75t_R register___U3690 ( .A(register__n2889), .Y(register__n3466) );
  AOI22xp33_ASAP7_75t_R register___U3691 ( .A1(register__n3393), .A2(register__n344), .B1(register__n1108), .B2(register__n337), 
        .Y(register__n12734) );
  CKINVDCx20_ASAP7_75t_R register___U3692 ( .A(register__n9750), .Y(register__n1108) );
  AND2x4_ASAP7_75t_R register___U3693 ( .A(RegWrite), .B(WB_rd[4]), .Y(register__n12483)
         );
  INVx1_ASAP7_75t_R register___U3694 ( .A(register__n13080), .Y(register__n1109) );
  BUFx3_ASAP7_75t_R register___U3695 ( .A(register__n5173), .Y(register__n3918) );
  INVx2_ASAP7_75t_R register___U3696 ( .A(register__n11733), .Y(register__n1312) );
  BUFx6f_ASAP7_75t_R register___U3697 ( .A(register__net117890), .Y(register__net117889) );
  AOI211x1_ASAP7_75t_R register___U3698 ( .A1(register__n924), .A2(register__net93456), .B(register__n2517), .C(register__n2519), 
        .Y(register__n2523) );
  BUFx12f_ASAP7_75t_R register___U3699 ( .A(register__net128430), .Y(register__net91921) );
  BUFx6f_ASAP7_75t_R register___U3700 ( .A(register__net145052), .Y(register__net145051) );
  BUFx6f_ASAP7_75t_R register___U3701 ( .A(register__net136188), .Y(register__net139025) );
  HB1xp67_ASAP7_75t_R register___U3702 ( .A(register__n2890), .Y(register__n2889) );
  INVxp67_ASAP7_75t_R register___U3703 ( .A(register__n11941), .Y(register__n11928) );
  BUFx6f_ASAP7_75t_R register___U3704 ( .A(register__n11947), .Y(register__n3535) );
  INVx2_ASAP7_75t_R register___U3705 ( .A(register__n11946), .Y(register__n11927) );
  AND2x2_ASAP7_75t_R register___U3706 ( .A(register__n11728), .B(register__n772), .Y(register__C6423_net61355) );
  BUFx2_ASAP7_75t_R register___U3707 ( .A(register__net62886), .Y(register__net124979) );
  HB1xp67_ASAP7_75t_R register___U3708 ( .A(register__n3431), .Y(register__n3430) );
  HB1xp67_ASAP7_75t_R register___U3709 ( .A(register__n3426), .Y(register__n4954) );
  CKINVDCx5p33_ASAP7_75t_R register___U3710 ( .A(register__net64976), .Y(register__net64940) );
  INVxp67_ASAP7_75t_R register___U3711 ( .A(register__n1794), .Y(register__n1617) );
  AO22x1_ASAP7_75t_R register___U3712 ( .A1(register__n9315), .A2(register__n481), .B1(register__n9417), .B2(register__n639), .Y(
        n11699) );
  AND3x2_ASAP7_75t_R register___U3713 ( .A(WB_rd[2]), .B(WB_rd[0]), .C(
        n5735), .Y(register__n12484) );
  HB1xp67_ASAP7_75t_R register___U3714 ( .A(register__n11655), .Y(register__n2890) );
  INVxp33_ASAP7_75t_R register___U3715 ( .A(register__n353), .Y(register__n1115) );
  INVxp33_ASAP7_75t_R register___U3716 ( .A(register__n353), .Y(register__n1116) );
  HB1xp67_ASAP7_75t_R register___U3717 ( .A(register__n13029), .Y(register__n3401) );
  BUFx12f_ASAP7_75t_R register___U3718 ( .A(register__net130079), .Y(register__C6423_net69182) );
  NOR2xp33_ASAP7_75t_R register___U3719 ( .A(register__n9674), .B(register__n6430), .Y(register__n8606) );
  INVxp67_ASAP7_75t_R register___U3720 ( .A(register__n5006), .Y(register__n7285) );
  HB1xp67_ASAP7_75t_R register___U3721 ( .A(register__n5007), .Y(register__n5006) );
  BUFx6f_ASAP7_75t_R register___U3722 ( .A(register__n4377), .Y(register__n11936) );
  BUFx6f_ASAP7_75t_R register___U3723 ( .A(register__net139925), .Y(register__net139924) );
  BUFx6f_ASAP7_75t_R register___U3724 ( .A(register__net62886), .Y(register__net139925) );
  INVx1_ASAP7_75t_R register___U3725 ( .A(register__n13070), .Y(register__n1119) );
  INVx1_ASAP7_75t_R register___U3726 ( .A(register__n13254), .Y(register__n1121) );
  AOI22xp5_ASAP7_75t_R register___U3727 ( .A1(register__net62864), .A2(register__n1726), .B1(register__n1122), .B2(
        n1699), .Y(register__n13241) );
  CKINVDCx20_ASAP7_75t_R register___U3728 ( .A(register__net89565), .Y(register__n1122) );
  INVx3_ASAP7_75t_R register___U3729 ( .A(register__net62864), .Y(register__net62820) );
  INVx1_ASAP7_75t_R register___U3730 ( .A(register__n13253), .Y(register__n1123) );
  NAND2xp67_ASAP7_75t_R register___U3731 ( .A(register__net91255), .B(register__n1115), .Y(register__n2583) );
  NAND2xp33_ASAP7_75t_R register___U3732 ( .A(register__n2015), .B(register__n2460), .Y(register__n2447) );
  INVxp67_ASAP7_75t_R register___U3733 ( .A(register__n3714), .Y(register__n5384) );
  HB1xp67_ASAP7_75t_R register___U3734 ( .A(register__n3715), .Y(register__n3714) );
  OAI22xp5_ASAP7_75t_R register___U3735 ( .A1(register__n4045), .A2(register__n1836), .B1(register__n6051), .B2(register__n1696), 
        .Y(register__n1125) );
  BUFx3_ASAP7_75t_R register___U3736 ( .A(register__net91921), .Y(register__net64964) );
  INVx1_ASAP7_75t_R register___U3737 ( .A(register__n2743), .Y(register__n1165) );
  BUFx5_ASAP7_75t_R register___U3738 ( .A(register__net62884), .Y(register__net62868) );
  AO22x1_ASAP7_75t_R register___U3739 ( .A1(register__n12330), .A2(register__n1721), .B1(register__n1127), .B2(register__n1712), 
        .Y(register__n1126) );
  CKINVDCx20_ASAP7_75t_R register___U3740 ( .A(register__n10003), .Y(register__n1127) );
  INVx3_ASAP7_75t_R register___U3741 ( .A(register__n12330), .Y(register__n12312) );
  BUFx6f_ASAP7_75t_R register___U3742 ( .A(register__n12500), .Y(register__n11809) );
  HB1xp67_ASAP7_75t_R register___U3743 ( .A(register__net63054), .Y(register__net145052) );
  HB1xp67_ASAP7_75t_R register___U3744 ( .A(register__n12983), .Y(register__n4155) );
  CKINVDCx20_ASAP7_75t_R register___U3745 ( .A(register__n9977), .Y(register__n1130) );
  HB1xp67_ASAP7_75t_R register___U3746 ( .A(register__n12721), .Y(register__n3787) );
  OAI22xp33_ASAP7_75t_R register___U3747 ( .A1(register__n12120), .A2(register__n2220), .B1(register__n10231), .B2(
        n11809), .Y(register__n2204) );
  HB1xp67_ASAP7_75t_R register___U3748 ( .A(register__n13325), .Y(register__n3715) );
  INVx1_ASAP7_75t_R register___U3749 ( .A(register__n12713), .Y(register__n1132) );
  INVxp67_ASAP7_75t_R register___U3750 ( .A(register__n4204), .Y(register__n7284) );
  HB1xp67_ASAP7_75t_R register___U3751 ( .A(register__n4205), .Y(register__n4204) );
  BUFx12f_ASAP7_75t_R register___U3752 ( .A(register__n2846), .Y(register__n11797) );
  AND2x2_ASAP7_75t_R register___U3753 ( .A(register__n1948), .B(register__n12485), .Y(register__n12486) );
  INVx6_ASAP7_75t_R register___U3754 ( .A(register__C6423_net69182), .Y(register__n_cell_125217_net175364) );
  HB1xp67_ASAP7_75t_R register___U3755 ( .A(register__n2843), .Y(register__n2136) );
  NOR2xp33_ASAP7_75t_R register___U3756 ( .A(register__C6422_net60224), .B(register__n1995), .Y(register__n2424) );
  HB1xp67_ASAP7_75t_R register___U3757 ( .A(register__n11198), .Y(register__n5332) );
  OAI22xp5_ASAP7_75t_R register___U3758 ( .A1(register__net66312), .A2(register__n6162), .B1(register__n5497), .B2(
        n1687), .Y(read_reg_data_2[20]) );
  AOI22xp33_ASAP7_75t_R register___U3759 ( .A1(register__n3729), .A2(register__n307), .B1(register__n1244), .B2(register__n4269), 
        .Y(register__n12693) );
  BUFx4f_ASAP7_75t_R register___U3760 ( .A(register__n3179), .Y(register__n3178) );
  HB1xp67_ASAP7_75t_R register___U3761 ( .A(register__n13211), .Y(register__n4530) );
  AO22x1_ASAP7_75t_R register___U3762 ( .A1(register__n9252), .A2(register__C6423_net61326), .B1(register__n10056), 
        .B2(register__C6423_net61325), .Y(register__n11528) );
  AO22x1_ASAP7_75t_R register___U3763 ( .A1(register__n9250), .A2(register__n1035), .B1(register__n7457), .B2(register__n2001), 
        .Y(register__n11549) );
  AO22x1_ASAP7_75t_R register___U3764 ( .A1(register__n9248), .A2(register__C6423_net68950), .B1(register__n10052), 
        .B2(register__n2000), .Y(register__n11568) );
  BUFx12f_ASAP7_75t_R register___U3765 ( .A(register__n748), .Y(register__n1136) );
  INVxp67_ASAP7_75t_R register___U3766 ( .A(register__net36445), .Y(register__n1152) );
  NOR2xp67_ASAP7_75t_R register___U3767 ( .A(register__n2305), .B(register__n1890), .Y(register__net36445) );
  INVxp33_ASAP7_75t_R register___U3768 ( .A(register__n12378), .Y(register__n1153) );
  INVxp33_ASAP7_75t_R register___U3769 ( .A(register__n3300), .Y(register__n12378) );
  NAND2xp33_ASAP7_75t_R register___U3770 ( .A(register__n1608), .B(register__n3343), .Y(register__n1155) );
  INVxp33_ASAP7_75t_R register___U3771 ( .A(register__n9913), .Y(register__n1608) );
  HB1xp67_ASAP7_75t_R register___U3772 ( .A(register__n12383), .Y(register__n3410) );
  INVxp67_ASAP7_75t_R register___U3773 ( .A(register__n6499), .Y(register__n7031) );
  HB1xp67_ASAP7_75t_R register___U3774 ( .A(register__n13084), .Y(register__n6499) );
  INVx1_ASAP7_75t_R register___U3775 ( .A(register__n12602), .Y(register__n1156) );
  AO22x1_ASAP7_75t_R register___U3776 ( .A1(register__n12295), .A2(register__n3354), .B1(register__n1158), .B2(register__n1711), 
        .Y(register__n1157) );
  CKINVDCx20_ASAP7_75t_R register___U3777 ( .A(register__n10243), .Y(register__n1158) );
  AND2x2_ASAP7_75t_R register___U3778 ( .A(register__net108812), .B(register__n1653), .Y(register__n2310) );
  HB1xp67_ASAP7_75t_R register___U3779 ( .A(register__C6423_net61194), .Y(register__net108812) );
  BUFx3_ASAP7_75t_R register___U3780 ( .A(register__n11419), .Y(register__n4910) );
  BUFx12f_ASAP7_75t_R register___U3781 ( .A(register__n3284), .Y(register__n3266) );
  INVxp67_ASAP7_75t_R register___U3782 ( .A(register__n3788), .Y(register__n5718) );
  BUFx3_ASAP7_75t_R register___U3783 ( .A(register__n10783), .Y(register__n5475) );
  INVx6_ASAP7_75t_R register___U3784 ( .A(register__net64464), .Y(register__net64430) );
  HB1xp67_ASAP7_75t_R register___U3785 ( .A(register__n4127), .Y(register__n1162) );
  HB1xp67_ASAP7_75t_R register___U3786 ( .A(register__n4127), .Y(register__n1163) );
  BUFx2_ASAP7_75t_R register___U3787 ( .A(register__n11730), .Y(register__n3719) );
  AO22x1_ASAP7_75t_R register___U3788 ( .A1(register__n7401), .A2(register__net146317), .B1(register__n5649), .B2(
        C6423_net74857), .Y(register__n1167) );
  AOI21x1_ASAP7_75t_R register___U3789 ( .A1(register__net125797), .A2(register__net93396), .B(register__n2497), .Y(
        n2516) );
  AO22x1_ASAP7_75t_R register___U3790 ( .A1(register__n8767), .A2(register__C6422_net70282), .B1(register__n9361), .B2(
        C6422_net70296), .Y(register__n10832) );
  BUFx12f_ASAP7_75t_R register___U3791 ( .A(register__n4633), .Y(register__n12126) );
  INVx1_ASAP7_75t_R register___U3792 ( .A(register__n11614), .Y(register__n1168) );
  INVxp67_ASAP7_75t_R register___U3793 ( .A(register__n1722), .Y(register__n1723) );
  INVxp67_ASAP7_75t_R register___U3794 ( .A(register__n1725), .Y(register__n1726) );
  INVxp67_ASAP7_75t_R register___U3795 ( .A(register__n1727), .Y(register__n1728) );
  INVx4_ASAP7_75t_R register___U3796 ( .A(register__n3353), .Y(register__n1738) );
  INVxp67_ASAP7_75t_R register___U3797 ( .A(register__n5413), .Y(register__n1575) );
  HB1xp67_ASAP7_75t_R register___U3798 ( .A(register__n6146), .Y(register__n5413) );
  AO22x1_ASAP7_75t_R register___U3799 ( .A1(register__n7809), .A2(register__net123861), .B1(register__n6878), .B2(
        C6423_net69198), .Y(register__n11421) );
  BUFx3_ASAP7_75t_R register___U3800 ( .A(register__net141083), .Y(register__net123861) );
  OA22x2_ASAP7_75t_R register___U3801 ( .A1(register__net62822), .A2(register__n1576), .B1(register__net89013), .B2(
        n2135), .Y(register__n12890) );
  BUFx3_ASAP7_75t_R register___U3802 ( .A(register__net103352), .Y(register__net89013) );
  INVxp67_ASAP7_75t_R register___U3803 ( .A(register__n6789), .Y(register__n7903) );
  BUFx3_ASAP7_75t_R register___U3804 ( .A(register__net129787), .Y(register__C6423_net69272) );
  BUFx3_ASAP7_75t_R register___U3805 ( .A(register__net128125), .Y(register__net101424) );
  BUFx6f_ASAP7_75t_R register___U3806 ( .A(register__net101424), .Y(register__C6423_net69250) );
  INVx2_ASAP7_75t_R register___U3807 ( .A(register__C6423_net69250), .Y(register__n_cell_124679_net156005) );
  OAI22xp5_ASAP7_75t_R register___U3808 ( .A1(register__net64440), .A2(register__n7327), .B1(register__net117709), .B2(
        n11834), .Y(register__n1250) );
  INVx6_ASAP7_75t_R register___U3809 ( .A(register__net64470), .Y(register__net64440) );
  INVxp67_ASAP7_75t_R register___U3810 ( .A(register__n4154), .Y(register__n5388) );
  HB1xp67_ASAP7_75t_R register___U3811 ( .A(register__n4155), .Y(register__n4154) );
  OAI22xp5_ASAP7_75t_R register___U3812 ( .A1(register__net64440), .A2(register__n113), .B1(register__net104579), .B2(
        n1528), .Y(register__n1253) );
  NOR2xp67_ASAP7_75t_R register___U3813 ( .A(register__n12172), .B(register__n1974), .Y(register__n1169) );
  NOR2xp33_ASAP7_75t_R register___U3814 ( .A(register__n1169), .B(register__n1170), .Y(register__n12904) );
  INVx1_ASAP7_75t_R register___U3815 ( .A(register__net36437), .Y(register__n1173) );
  INVx1_ASAP7_75t_R register___U3816 ( .A(register__n13322), .Y(register__n1174) );
  INVxp67_ASAP7_75t_R register___U3817 ( .A(register__n12979), .Y(register__n3751) );
  AO21x1_ASAP7_75t_R register___U3818 ( .A1(register__n128), .A2(register__net90217), .B(register__n1175), .Y(register__n2578) );
  AND2x2_ASAP7_75t_R register___U3819 ( .A(register__net125170), .B(register__net90229), .Y(register__n1175) );
  BUFx6f_ASAP7_75t_R register___U3820 ( .A(register__n3354), .Y(register__n3352) );
  BUFx6f_ASAP7_75t_R register___U3821 ( .A(register__n3298), .Y(register__n3564) );
  BUFx6f_ASAP7_75t_R register___U3822 ( .A(register__n6269), .Y(register__n12440) );
  BUFx12f_ASAP7_75t_R register___U3823 ( .A(register__n11739), .Y(register__n3075) );
  INVxp67_ASAP7_75t_R register___U3824 ( .A(register__n12914), .Y(register__n4385) );
  AO22x1_ASAP7_75t_R register___U3825 ( .A1(register__net88584), .A2(register__n1853), .B1(register__net88500), .B2(
        net139537), .Y(register__n10811) );
  HB1xp67_ASAP7_75t_R register___U3826 ( .A(register__n13009), .Y(register__n3890) );
  HB1xp67_ASAP7_75t_R register___U3827 ( .A(register__n6790), .Y(register__n6789) );
  BUFx6f_ASAP7_75t_R register___U3828 ( .A(register__net124977), .Y(register__net140665) );
  INVx2_ASAP7_75t_R register___U3829 ( .A(register__n5739), .Y(register__n8255) );
  INVx1_ASAP7_75t_R register___U3830 ( .A(register__n1736), .Y(register__n1737) );
  INVx1_ASAP7_75t_R register___U3831 ( .A(register__n13238), .Y(register__n1176) );
  NOR2x2_ASAP7_75t_R register___U3832 ( .A(register__n4582), .B(register__n1178), .Y(register__n1177) );
  INVx3_ASAP7_75t_R register___U3833 ( .A(register__n12444), .Y(register__n12422) );
  INVxp67_ASAP7_75t_R register___U3834 ( .A(register__n3889), .Y(register__n8603) );
  HB1xp67_ASAP7_75t_R register___U3835 ( .A(register__n3890), .Y(register__n3889) );
  AO22x1_ASAP7_75t_R register___U3836 ( .A1(register__n9842), .A2(register__net93569), .B1(register__n10267), .B2(register__n284), 
        .Y(register__n11655) );
  OA22x2_ASAP7_75t_R register___U3837 ( .A1(register__n12426), .A2(register__n335), .B1(register__n9895), .B2(register__n68), .Y(
        n12720) );
  HB1xp67_ASAP7_75t_R register___U3838 ( .A(register__n3840), .Y(register__n6266) );
  INVxp33_ASAP7_75t_R register___U3839 ( .A(register__net125170), .Y(register__n1179) );
  INVx2_ASAP7_75t_R register___U3840 ( .A(register__net125169), .Y(register__n1180) );
  INVx2_ASAP7_75t_R register___U3841 ( .A(register__net125169), .Y(register__n1181) );
  AND2x2_ASAP7_75t_R register___U3842 ( .A(register__n11279), .B(register__n11278), .Y(register__n1182) );
  AND3x1_ASAP7_75t_R register___U3843 ( .A(register__n1182), .B(register__n9232), .C(register__n11280), .Y(register__n8640) );
  BUFx2_ASAP7_75t_R register___U3844 ( .A(register__net125170), .Y(register__net125169) );
  OAI22xp5_ASAP7_75t_R register___U3845 ( .A1(register__net66304), .A2(register__n8640), .B1(register__net64780), .B2(
        n1687), .Y(read_reg_data_2[6]) );
  BUFx6f_ASAP7_75t_R register___U3846 ( .A(register__net139924), .Y(register__net62860) );
  INVx1_ASAP7_75t_R register___U3847 ( .A(register__n1567), .Y(register__n1183) );
  INVx1_ASAP7_75t_R register___U3848 ( .A(register__n118), .Y(register__register__n1184) );
  INVxp67_ASAP7_75t_R register___U3849 ( .A(register__n1922), .Y(register__n1185) );
  INVxp67_ASAP7_75t_R register___U3850 ( .A(register__n118), .Y(register__register__n1186) );
  INVx1_ASAP7_75t_R register___U3851 ( .A(register__n1566), .Y(register__n1187) );
  INVxp33_ASAP7_75t_R register___U3852 ( .A(register__n1564), .Y(register__n1188) );
  INVxp67_ASAP7_75t_R register___U3853 ( .A(register__n1922), .Y(register__n1189) );
  INVxp67_ASAP7_75t_R register___U3854 ( .A(register__n1565), .Y(register__n1190) );
  INVxp67_ASAP7_75t_R register___U3855 ( .A(register__n2140), .Y(register__n1191) );
  INVxp67_ASAP7_75t_R register___U3856 ( .A(register__n1922), .Y(register__n1192) );
  INVxp33_ASAP7_75t_R register___U3857 ( .A(register__n1568), .Y(register__n1193) );
  INVx1_ASAP7_75t_R register___U3858 ( .A(register__n1569), .Y(register__n1195) );
  INVx1_ASAP7_75t_R register___U3859 ( .A(register__n1568), .Y(register__n1196) );
  INVx1_ASAP7_75t_R register___U3860 ( .A(register__n1567), .Y(register__n1197) );
  INVx1_ASAP7_75t_R register___U3861 ( .A(register__n1565), .Y(register__n1198) );
  INVx1_ASAP7_75t_R register___U3862 ( .A(register__n1564), .Y(register__n1199) );
  INVx1_ASAP7_75t_R register___U3863 ( .A(register__n1566), .Y(register__n1200) );
  INVxp33_ASAP7_75t_R register___U3864 ( .A(register__net74029), .Y(register__n1201) );
  INVxp67_ASAP7_75t_R register___U3865 ( .A(register__n2144), .Y(register__n1202) );
  INVxp67_ASAP7_75t_R register___U3866 ( .A(register__n2150), .Y(register__n1205) );
  INVx2_ASAP7_75t_R register___U3867 ( .A(register__n2146), .Y(register__n1206) );
  INVx1_ASAP7_75t_R register___U3868 ( .A(register__n2152), .Y(register__n1207) );
  INVx1_ASAP7_75t_R register___U3869 ( .A(register__net67382), .Y(register__n1208) );
  INVx1_ASAP7_75t_R register___U3870 ( .A(register__n2154), .Y(register__n1209) );
  INVx1_ASAP7_75t_R register___U3871 ( .A(register__n2148), .Y(register__n1210) );
  INVx6_ASAP7_75t_R register___U3872 ( .A(register__net74013), .Y(register__n1212) );
  INVxp67_ASAP7_75t_R register___U3873 ( .A(register__n1563), .Y(register__n1564) );
  INVx2_ASAP7_75t_R register___U3874 ( .A(register__n2145), .Y(register__n2146) );
  INVx1_ASAP7_75t_R register___U3875 ( .A(register__n2153), .Y(register__n2154) );
  INVxp33_ASAP7_75t_R register___U3876 ( .A(register__net106927), .Y(register__n2142) );
  BUFx12f_ASAP7_75t_R register___U3877 ( .A(register__n1194), .Y(register__net67414) );
  INVx1_ASAP7_75t_R register___U3878 ( .A(register__net74029), .Y(register__net73977) );
  INVx1_ASAP7_75t_R register___U3879 ( .A(register__net67382), .Y(register__n2153) );
  INVx1_ASAP7_75t_R register___U3880 ( .A(register__n13102), .Y(register__n1213) );
  BUFx3_ASAP7_75t_R register___U3881 ( .A(register__net141041), .Y(register__net141039) );
  HB1xp67_ASAP7_75t_R register___U3882 ( .A(register__n12553), .Y(register__n6251) );
  BUFx6f_ASAP7_75t_R register___U3883 ( .A(register__net143517), .Y(register__net143790) );
  BUFx2_ASAP7_75t_R register___U3884 ( .A(register__n4583), .Y(register__n4582) );
  HB1xp67_ASAP7_75t_R register___U3885 ( .A(register__n11331), .Y(register__n4583) );
  INVx2_ASAP7_75t_R register___U3886 ( .A(register__n1483), .Y(register__n1484) );
  NOR2x2_ASAP7_75t_R register___U3887 ( .A(register__n5302), .B(register__n4625), .Y(register__n1483) );
  INVx2_ASAP7_75t_R register___U3888 ( .A(register__n3308), .Y(register__n1790) );
  INVxp67_ASAP7_75t_R register___U3889 ( .A(register__n5779), .Y(register__n8665) );
  INVx1_ASAP7_75t_R register___U3890 ( .A(register__n2306), .Y(register__n1890) );
  AO22x1_ASAP7_75t_R register___U3891 ( .A1(register__n6943), .A2(register__C6423_net61318), .B1(register__n10241), 
        .B2(register__n1451), .Y(register__n11507) );
  AO22x1_ASAP7_75t_R register___U3892 ( .A1(register__n9814), .A2(register__C6423_net61318), .B1(register__n8157), .B2(
        n1453), .Y(register__n11376) );
  AO22x1_ASAP7_75t_R register___U3893 ( .A1(register__n7549), .A2(register__n128), .B1(register__n7841), .B2(register__n1449), 
        .Y(register__n11712) );
  INVxp67_ASAP7_75t_R register___U3894 ( .A(register__net124439), .Y(register__net109491) );
  AO22x1_ASAP7_75t_R register___U3895 ( .A1(register__n9905), .A2(register__net137440), .B1(register__n6385), .B2(
        net139058), .Y(register__n11419) );
  BUFx2_ASAP7_75t_R register___U3896 ( .A(register__n7351), .Y(register__n7350) );
  NAND2xp33_ASAP7_75t_R register___U3897 ( .A(register__n10491), .B(register__net125170), .Y(register__n1214) );
  NAND2xp33_ASAP7_75t_R register___U3898 ( .A(register__n8785), .B(register__net94399), .Y(register__n1215) );
  NAND2xp67_ASAP7_75t_R register___U3899 ( .A(register__n1214), .B(register__n1215), .Y(register__n11330) );
  INVx2_ASAP7_75t_R register___U3900 ( .A(register__n11330), .Y(register__n8277) );
  INVxp67_ASAP7_75t_R register___U3901 ( .A(register__n5407), .Y(register__n6688) );
  HB1xp67_ASAP7_75t_R register___U3902 ( .A(register__n5408), .Y(register__n5407) );
  NOR3xp33_ASAP7_75t_R register___U3903 ( .A(register__n1562), .B(register__n1289), .C(register__n11618), .Y(register__n1216) );
  NOR2xp67_ASAP7_75t_R register___U3904 ( .A(register__n1561), .B(register__n1217), .Y(register__n8585) );
  INVxp67_ASAP7_75t_R register___U3905 ( .A(register__n1216), .Y(register__n1217) );
  INVx1_ASAP7_75t_R register___U3906 ( .A(register__n11617), .Y(register__n1561) );
  NAND4xp25_ASAP7_75t_R register___U3907 ( .A(register__n1472), .B(register__n5702), .C(register__n8229), .D(register__n2259), 
        .Y(register__n1562) );
  OAI21xp33_ASAP7_75t_R register___U3908 ( .A1(register__n420), .A2(register__n2638), .B(register__n2664), .Y(register__n2665) );
  INVx1_ASAP7_75t_R register___U3909 ( .A(register__n13109), .Y(register__n1218) );
  BUFx3_ASAP7_75t_R register___U3910 ( .A(register__n4929), .Y(register__n4928) );
  HB1xp67_ASAP7_75t_R register___U3911 ( .A(register__n12922), .Y(register__n3957) );
  HB1xp67_ASAP7_75t_R register___U3912 ( .A(register__n13342), .Y(register__n7351) );
  INVx1_ASAP7_75t_R register___U3913 ( .A(register__n3754), .Y(register__n12320) );
  NOR2xp67_ASAP7_75t_R register___U3914 ( .A(register__n1219), .B(register__n1220), .Y(register__n7274) );
  NAND2xp67_ASAP7_75t_R register___U3915 ( .A(register__n11561), .B(register__n11562), .Y(register__n1219) );
  NAND2xp67_ASAP7_75t_R register___U3916 ( .A(register__n11560), .B(register__n7959), .Y(register__n1220) );
  INVx1_ASAP7_75t_R register___U3917 ( .A(register__n12326), .Y(register__n12313) );
  HB1xp67_ASAP7_75t_R register___U3918 ( .A(register__n3789), .Y(register__n3788) );
  OAI21xp33_ASAP7_75t_R register___U3919 ( .A1(register__C6423_net68516), .A2(register__n2532), .B(register__n2563), 
        .Y(register__n2562) );
  INVxp67_ASAP7_75t_R register___U3920 ( .A(register__n3769), .Y(register__n6184) );
  HB1xp67_ASAP7_75t_R register___U3921 ( .A(register__n13288), .Y(register__n4674) );
  INVx1_ASAP7_75t_R register___U3922 ( .A(register__n13309), .Y(register__n1221) );
  INVx1_ASAP7_75t_R register___U3923 ( .A(register__n11171), .Y(register__n1222) );
  BUFx2_ASAP7_75t_R register___U3924 ( .A(register__n10525), .Y(register__n5125) );
  INVxp67_ASAP7_75t_R register___U3925 ( .A(register__n10528), .Y(register__n8303) );
  INVxp67_ASAP7_75t_R register___U3926 ( .A(register__n4673), .Y(register__n6696) );
  HB1xp67_ASAP7_75t_R register___U3927 ( .A(register__n4674), .Y(register__n4673) );
  AND4x2_ASAP7_75t_R register___U3928 ( .A(register__n6701), .B(register__n1505), .C(register__n6700), .D(register__n5252), .Y(
        n11155) );
  INVx2_ASAP7_75t_R register___U3929 ( .A(register__n11166), .Y(register__n6701) );
  INVx1_ASAP7_75t_R register___U3930 ( .A(register__n12728), .Y(register__n1223) );
  AOI22xp33_ASAP7_75t_R register___U3931 ( .A1(register__net138885), .A2(register__n1379), .B1(register__n1380), .B2(
        n1381), .Y(register__n12838) );
  INVx1_ASAP7_75t_R register___U3932 ( .A(register__n11309), .Y(register__n1224) );
  HB1xp67_ASAP7_75t_R register___U3933 ( .A(register__n5780), .Y(register__n5779) );
  HB1xp67_ASAP7_75t_R register___U3934 ( .A(register__n13101), .Y(register__n5780) );
  HB1xp67_ASAP7_75t_R register___U3935 ( .A(register__n12814), .Y(register__n5408) );
  BUFx3_ASAP7_75t_R register___U3936 ( .A(register__n12932), .Y(register__n3977) );
  AOI22xp33_ASAP7_75t_R register___U3937 ( .A1(register__net90261), .A2(register__C6423_net61343), .B1(
        net89421), .B2(register__net122313), .Y(register__n1407) );
  HB1xp67_ASAP7_75t_R register___U3938 ( .A(register__n13074), .Y(register__n4676) );
  HB1xp67_ASAP7_75t_R register___U3939 ( .A(register__n3770), .Y(register__n3769) );
  BUFx6f_ASAP7_75t_R register___U3940 ( .A(register__net64818), .Y(register__net105198) );
  INVx2_ASAP7_75t_R register___U3941 ( .A(register__n1793), .Y(register__n1642) );
  HB1xp67_ASAP7_75t_R register___U3942 ( .A(register__n4776), .Y(register__n4775) );
  INVx1_ASAP7_75t_R register___U3943 ( .A(register__n13150), .Y(register__n1227) );
  HB1xp67_ASAP7_75t_R register___U3944 ( .A(register__net63390), .Y(register__net141997) );
  BUFx6f_ASAP7_75t_R register___U3945 ( .A(register__net64380), .Y(register__net64392) );
  INVxp67_ASAP7_75t_R register___U3946 ( .A(register__n3786), .Y(register__n8594) );
  HB1xp67_ASAP7_75t_R register___U3947 ( .A(register__n3787), .Y(register__n3786) );
  HB1xp67_ASAP7_75t_R register___U3948 ( .A(register__n13323), .Y(register__n3789) );
  CKINVDCx20_ASAP7_75t_R register___U3949 ( .A(register__n1570), .Y(register__n1228) );
  AO22x1_ASAP7_75t_R register___U3950 ( .A1(register__n9704), .A2(register__n85), .B1(register__n10034), .B2(register__n422), .Y(
        n11555) );
  AO22x1_ASAP7_75t_R register___U3951 ( .A1(register__n9670), .A2(register__net150060), .B1(register__n9917), .B2(register__n2024), .Y(register__n11556) );
  BUFx3_ASAP7_75t_R register___U3952 ( .A(register__n3977), .Y(register__n3976) );
  OAI22xp5_ASAP7_75t_R register___U3953 ( .A1(register__net66314), .A2(register__n7274), .B1(register__n3410), .B2(
        n1687), .Y(read_reg_data_2[22]) );
  AND2x2_ASAP7_75t_R register___U3954 ( .A(register__n7930), .B(register__n1555), .Y(register__n1229) );
  HB1xp67_ASAP7_75t_R register___U3955 ( .A(register__n4635), .Y(register__n12129) );
  AO22x1_ASAP7_75t_R register___U3956 ( .A1(register__n9680), .A2(register__net109204), .B1(register__n9927), .B2(
        net129911), .Y(register__n10542) );
  NOR2xp33_ASAP7_75t_R register___U3957 ( .A(register__n1172), .B(register__n2593), .Y(register__n2595) );
  INVx1_ASAP7_75t_R register___U3958 ( .A(register__n12778), .Y(register__n1231) );
  AOI22xp33_ASAP7_75t_R register___U3959 ( .A1(register__net62874), .A2(register__n3336), .B1(register__n2543), .B2(
        n1755), .Y(register__n13118) );
  HB1xp67_ASAP7_75t_R register___U3960 ( .A(register__net124977), .Y(register__net62874) );
  NOR2xp33_ASAP7_75t_R register___U3961 ( .A(register__n1232), .B(register__n1233), .Y(register__n1234) );
  NOR2xp67_ASAP7_75t_R register___U3962 ( .A(register__n1234), .B(register__n2581), .Y(register__n2527) );
  INVxp33_ASAP7_75t_R register___U3963 ( .A(register__net93661), .Y(register__n1232) );
  INVxp33_ASAP7_75t_R register___U3964 ( .A(register__n1452), .Y(register__n1233) );
  BUFx3_ASAP7_75t_R register___U3965 ( .A(register__net101126), .Y(register__net93661) );
  INVx1_ASAP7_75t_R register___U3966 ( .A(register__n12951), .Y(register__n1235) );
  AND3x2_ASAP7_75t_R register___U3967 ( .A(register__n1513), .B(register__n11143), .C(register__n11132), .Y(register__n11141) );
  INVx1_ASAP7_75t_R register___U3968 ( .A(register__n12981), .Y(register__n1236) );
  INVx1_ASAP7_75t_R register___U3969 ( .A(register__n11193), .Y(register__n1237) );
  INVx1_ASAP7_75t_R register___U3970 ( .A(register__n11121), .Y(register__n1260) );
  AND4x2_ASAP7_75t_R register___U3971 ( .A(register__n1611), .B(register__n3345), .C(register__n2225), .D(register__n3063), .Y(
        n11121) );
  AOI22xp33_ASAP7_75t_R register___U3972 ( .A1(register__net62874), .A2(register__n972), .B1(register__n2553), .B2(register__n979), .Y(register__n13179) );
  INVxp67_ASAP7_75t_R register___U3973 ( .A(register__n5167), .Y(register__n8325) );
  AO22x1_ASAP7_75t_R register___U3974 ( .A1(register__n9619), .A2(register__C6423_net61343), .B1(register__n10066), 
        .B2(register__net129787), .Y(register__n11166) );
  AO22x1_ASAP7_75t_R register___U3975 ( .A1(register__n10485), .A2(register__C6423_net61343), .B1(register__n10458), 
        .B2(register__net129787), .Y(register__n11188) );
  BUFx4f_ASAP7_75t_R register___U3976 ( .A(register__net125327), .Y(register__net129615) );
  OAI22xp5_ASAP7_75t_R register___U3977 ( .A1(register__net112762), .A2(register__n8338), .B1(register__n11965), .B2(
        n1687), .Y(read_reg_data_2[1]) );
  AO22x1_ASAP7_75t_R register___U3978 ( .A1(register__n9262), .A2(register__C6423_net61343), .B1(register__n10102), 
        .B2(register__net129787), .Y(register__n11398) );
  AO22x1_ASAP7_75t_R register___U3979 ( .A1(register__n9617), .A2(register__C6423_net61343), .B1(register__n8946), .B2(
        net129787), .Y(register__n11211) );
  AO22x1_ASAP7_75t_R register___U3980 ( .A1(register__n9812), .A2(register__C6423_net61343), .B1(register__n10142), 
        .B2(register__net129787), .Y(register__n11378) );
  BUFx6f_ASAP7_75t_R register___U3981 ( .A(register__n6267), .Y(register__n12438) );
  INVx2_ASAP7_75t_R register___U3982 ( .A(register__n4736), .Y(register__n8265) );
  NOR3xp33_ASAP7_75t_R register___U3983 ( .A(register__n2491), .B(register__n2486), .C(register__n2485), .Y(register__n1239) );
  NOR2xp33_ASAP7_75t_R register___U3984 ( .A(register__n2508), .B(register__n1240), .Y(register__n2507) );
  NOR2xp33_ASAP7_75t_R register___U3985 ( .A(register__n1172), .B(register__n2483), .Y(register__n2485) );
  NOR2x1p5_ASAP7_75t_R register___U3986 ( .A(register__n2484), .B(register__n1441), .Y(register__n2486) );
  INVx6_ASAP7_75t_R register___U3987 ( .A(register__net130020), .Y(register__net63258) );
  INVx1_ASAP7_75t_R register___U3988 ( .A(register__n13257), .Y(register__n1241) );
  BUFx6f_ASAP7_75t_R register___U3989 ( .A(write_data[7]), .Y(register__net64734) );
  INVx1_ASAP7_75t_R register___U3990 ( .A(register__n11358), .Y(register__n1242) );
  AOI21xp5_ASAP7_75t_R register___U3991 ( .A1(register__net139058), .A2(register__net89017), .B(register__n2578), .Y(
        n2579) );
  BUFx2_ASAP7_75t_R register___U3992 ( .A(register__n11691), .Y(register__n4622) );
  BUFx6f_ASAP7_75t_R register___U3993 ( .A(register__net124979), .Y(register__net62884) );
  BUFx3_ASAP7_75t_R register___U3994 ( .A(register__n11530), .Y(register__n5309) );
  HB1xp67_ASAP7_75t_R register___U3995 ( .A(register__net124979), .Y(register__net62872) );
  BUFx2_ASAP7_75t_R register___U3996 ( .A(register__n3077), .Y(register__n3371) );
  HB1xp67_ASAP7_75t_R register___U3997 ( .A(register__n3078), .Y(register__n3077) );
  HB1xp67_ASAP7_75t_R register___U3998 ( .A(register__n1084), .Y(register__n4913) );
  BUFx3_ASAP7_75t_R register___U3999 ( .A(register__net64720), .Y(register__net137456) );
  HB1xp67_ASAP7_75t_R register___U4000 ( .A(register__net144804), .Y(register__net64720) );
  BUFx3_ASAP7_75t_R register___U4001 ( .A(register__net144804), .Y(register__net64710) );
  INVxp67_ASAP7_75t_R register___U4002 ( .A(register__n4753), .Y(register__n8696) );
  HB1xp67_ASAP7_75t_R register___U4003 ( .A(register__n12629), .Y(register__n4416) );
  INVx1_ASAP7_75t_R register___U4004 ( .A(register__n10795), .Y(register__n1245) );
  INVx1_ASAP7_75t_R register___U4005 ( .A(register__n11275), .Y(register__n1246) );
  INVx6_ASAP7_75t_R register___U4006 ( .A(register__n12435), .Y(register__n7258) );
  AO22x1_ASAP7_75t_R register___U4007 ( .A1(register__n9601), .A2(register__n128), .B1(register__n10024), .B2(register__n1452), 
        .Y(register__n11331) );
  AO22x1_ASAP7_75t_R register___U4008 ( .A1(register__n9662), .A2(register__net125426), .B1(register__n9991), .B2(
        C6423_net68766), .Y(register__n11531) );
  BUFx3_ASAP7_75t_R register___U4009 ( .A(register__net120789), .Y(register__net120788) );
  AO22x1_ASAP7_75t_R register___U4010 ( .A1(register__n12385), .A2(register__n11752), .B1(register__n1488), .B2(register__n2834), 
        .Y(register__n1487) );
  INVxp67_ASAP7_75t_R register___U4011 ( .A(register__n7064), .Y(register__n4729) );
  NAND2xp67_ASAP7_75t_R register___U4012 ( .A(register__n1387), .B(register__n1386), .Y(register__n1554) );
  INVxp67_ASAP7_75t_R register___U4013 ( .A(register__net63290), .Y(register__n1552) );
  BUFx6f_ASAP7_75t_R register___U4014 ( .A(register__net124977), .Y(register__net62850) );
  NAND2xp67_ASAP7_75t_R register___U4015 ( .A(register__n1276), .B(register__n1277), .Y(register__n11592) );
  INVx1_ASAP7_75t_R register___U4016 ( .A(register__n12870), .Y(register__n1252) );
  BUFx6f_ASAP7_75t_R register___U4017 ( .A(register__n4746), .Y(register__n12302) );
  INVx1_ASAP7_75t_R register___U4018 ( .A(register__n12667), .Y(register__n1254) );
  AND2x2_ASAP7_75t_R register___U4019 ( .A(register__n1031), .B(register__n11298), .Y(register__n1255) );
  AND3x1_ASAP7_75t_R register___U4020 ( .A(register__n1255), .B(register__n11297), .C(register__n11299), .Y(register__n7613) );
  INVx6_ASAP7_75t_R register___U4021 ( .A(register__net129770), .Y(register__net129768) );
  BUFx12f_ASAP7_75t_R register___U4022 ( .A(register__net142360), .Y(register__net97625) );
  HB1xp67_ASAP7_75t_R register___U4023 ( .A(register__n4754), .Y(register__n4753) );
  HB1xp67_ASAP7_75t_R register___U4024 ( .A(register__n10592), .Y(register__n4754) );
  AO22x1_ASAP7_75t_R register___U4025 ( .A1(register__n8767), .A2(register__C6423_net61340), .B1(register__n9361), .B2(
        C6423_net69198), .Y(register__n11441) );
  AO22x1_ASAP7_75t_R register___U4026 ( .A1(register__n9847), .A2(register__C6423_net61340), .B1(register__n10167), 
        .B2(register__C6423_net69198), .Y(register__n11359) );
  INVx1_ASAP7_75t_R register___U4027 ( .A(register__n10852), .Y(register__n1256) );
  HB1xp67_ASAP7_75t_R register___U4028 ( .A(register__n4358), .Y(register__n4357) );
  AOI22xp33_ASAP7_75t_R register___U4029 ( .A1(register__net141489), .A2(register__n903), .B1(register__n1430), .B2(
        n891), .Y(register__n13058) );
  INVx1_ASAP7_75t_R register___U4030 ( .A(register__n12742), .Y(register__n1257) );
  BUFx6f_ASAP7_75t_R register___U4031 ( .A(register__n7592), .Y(register__n12417) );
  BUFx12f_ASAP7_75t_R register___U4032 ( .A(register__n12447), .Y(register__n3483) );
  INVx1_ASAP7_75t_R register___U4033 ( .A(register__n10565), .Y(register__n1258) );
  AND2x2_ASAP7_75t_R register___U4034 ( .A(register__n1258), .B(register__n1259), .Y(register__n10547) );
  INVx1_ASAP7_75t_R register___U4035 ( .A(register__n4377), .Y(register__n11921) );
  BUFx3_ASAP7_75t_R register___U4036 ( .A(register__n10780), .Y(register__n6705) );
  NAND3x1_ASAP7_75t_R register___U4037 ( .A(register__n1850), .B(register__n8249), .C(register__n8248), .Y(register__n1261) );
  AO22x1_ASAP7_75t_R register___U4038 ( .A1(register__n12268), .A2(register__n6160), .B1(register__n1264), .B2(register__n1703), 
        .Y(register__n1263) );
  NAND2x1p5_ASAP7_75t_R register___U4039 ( .A(register__n10268), .B(register__C6423_net69272), .Y(register__n1277) );
  INVxp67_ASAP7_75t_R register___U4040 ( .A(register__n5026), .Y(register__n7019) );
  AOI22xp33_ASAP7_75t_R register___U4041 ( .A1(register__n9630), .A2(register__n38), .B1(register__n10093), .B2(register__n369), 
        .Y(register__n1267) );
  CKINVDCx20_ASAP7_75t_R register___U4042 ( .A(register__net116000), .Y(register__n1269) );
  INVx2_ASAP7_75t_R register___U4043 ( .A(register__net64048), .Y(register__net64014) );
  HB1xp67_ASAP7_75t_R register___U4044 ( .A(register__n11670), .Y(register__n4358) );
  HB1xp67_ASAP7_75t_R register___U4045 ( .A(register__n13014), .Y(register__n3559) );
  INVxp67_ASAP7_75t_R register___U4046 ( .A(register__n3906), .Y(register__n5909) );
  HB1xp67_ASAP7_75t_R register___U4047 ( .A(register__n3907), .Y(register__n3906) );
  INVxp67_ASAP7_75t_R register___U4048 ( .A(register__n4423), .Y(register__n6686) );
  HB1xp67_ASAP7_75t_R register___U4049 ( .A(register__n4424), .Y(register__n4423) );
  INVxp67_ASAP7_75t_R register___U4050 ( .A(register__n3903), .Y(register__n4482) );
  INVx1_ASAP7_75t_R register___U4051 ( .A(register__n11099), .Y(register__n1271) );
  HB1xp67_ASAP7_75t_R register___U4052 ( .A(register__n12923), .Y(register__n3770) );
  INVx6_ASAP7_75t_R register___U4053 ( .A(register__net64916), .Y(register__net131433) );
  INVx1_ASAP7_75t_R register___U4054 ( .A(register__n11362), .Y(register__n1272) );
  BUFx6f_ASAP7_75t_R register___U4055 ( .A(register__net62886), .Y(register__net124977) );
  INVx6_ASAP7_75t_R register___U4056 ( .A(n11), .Y(register__net62886) );
  INVx1_ASAP7_75t_R register___U4057 ( .A(register__n13306), .Y(register__n1273) );
  HB1xp67_ASAP7_75t_R register___U4058 ( .A(register__n3421), .Y(register__n3754) );
  NAND3xp33_ASAP7_75t_R register___U4059 ( .A(register__n5704), .B(register__n5706), .C(register__n5705), .Y(register__n1274) );
  AOI22xp33_ASAP7_75t_R register___U4060 ( .A1(register__net64718), .A2(register__n1617), .B1(register__n1275), .B2(
        n1794), .Y(register__n12769) );
  CKINVDCx20_ASAP7_75t_R register___U4061 ( .A(register__n5681), .Y(register__n1275) );
  CKINVDCx5p33_ASAP7_75t_R register___U4062 ( .A(register__net64718), .Y(register__net64686) );
  BUFx2_ASAP7_75t_R register___U4063 ( .A(register__net140684), .Y(register__net145200) );
  BUFx3_ASAP7_75t_R register___U4064 ( .A(register__net140684), .Y(register__net145449) );
  BUFx3_ASAP7_75t_R register___U4065 ( .A(register__net140684), .Y(register__net63194) );
  NAND2x1_ASAP7_75t_R register___U4066 ( .A(register__n11658), .B(register__n6719), .Y(register__n2261) );
  AND4x2_ASAP7_75t_R register___U4067 ( .A(register__n6423), .B(register__n6422), .C(register__n5662), .D(register__n4355), .Y(
        n11658) );
  BUFx2_ASAP7_75t_R register___U4068 ( .A(register__n5031), .Y(register__n5030) );
  HB1xp67_ASAP7_75t_R register___U4069 ( .A(register__n12946), .Y(register__n4776) );
  BUFx12f_ASAP7_75t_R register___U4070 ( .A(register__net146677), .Y(register__net147289) );
  BUFx4f_ASAP7_75t_R register___U4071 ( .A(register__net91738), .Y(register__net140685) );
  INVx1_ASAP7_75t_R register___U4072 ( .A(register__n13153), .Y(register__n6440) );
  BUFx6f_ASAP7_75t_R register___U4073 ( .A(register__n8619), .Y(register__n3374) );
  BUFx6f_ASAP7_75t_R register___U4074 ( .A(register__n12417), .Y(register__n12409) );
  NAND2xp33_ASAP7_75t_R register___U4075 ( .A(register__n8769), .B(register__C6423_net61343), .Y(register__n1276) );
  OAI21xp33_ASAP7_75t_R register___U4076 ( .A1(register__n2489), .A2(register__n_cell_125217_net175396), .B(
        n2509), .Y(register__n2508) );
  NAND2xp33_ASAP7_75t_R register___U4077 ( .A(register__n2506), .B(register__n2507), .Y(register__n2464) );
  OAI21xp33_ASAP7_75t_R register___U4078 ( .A1(register__net66306), .A2(register__n2463), .B(register__n2467), .Y(
        read_reg_data_2[10]) );
  NOR2xp33_ASAP7_75t_R register___U4079 ( .A(register__net63342), .B(register__n335), .Y(register__n1279) );
  NOR2xp67_ASAP7_75t_R register___U4080 ( .A(register__n9830), .B(register__n345), .Y(register__n1280) );
  NOR2xp33_ASAP7_75t_R register___U4081 ( .A(register__n1279), .B(register__n1280), .Y(register__n12724) );
  INVx2_ASAP7_75t_R register___U4082 ( .A(register__net63366), .Y(register__net63334) );
  INVxp33_ASAP7_75t_R register___U4083 ( .A(register__net63376), .Y(register__net63342) );
  BUFx6f_ASAP7_75t_R register___U4084 ( .A(register__n7210), .Y(register__n9830) );
  NOR2xp67_ASAP7_75t_R register___U4085 ( .A(register__n2244), .B(register__n2245), .Y(register__n1303) );
  AO22x1_ASAP7_75t_R register___U4086 ( .A1(register__n9786), .A2(register__net125170), .B1(register__n10185), .B2(
        net94399), .Y(register__n11309) );
  HB1xp67_ASAP7_75t_R register___U4087 ( .A(register__n12669), .Y(register__n6784) );
  AO21x1_ASAP7_75t_R register___U4088 ( .A1(register__net89713), .A2(register__C6422_net70388), .B(register__n2340), 
        .Y(register__n2362) );
  BUFx2_ASAP7_75t_R register___U4089 ( .A(register__net123879), .Y(register__C6422_net70388) );
  AOI21x1_ASAP7_75t_R register___U4090 ( .A1(register__net126316), .A2(register__net90997), .B(register__n2362), .Y(
        n2361) );
  HB1xp67_ASAP7_75t_R register___U4091 ( .A(register__n10752), .Y(register__n5031) );
  INVxp67_ASAP7_75t_R register___U4092 ( .A(register__C6423_net69560), .Y(register__n2437) );
  INVx3_ASAP7_75t_R register___U4093 ( .A(register__n8226), .Y(register__n1480) );
  INVx3_ASAP7_75t_R register___U4094 ( .A(register__n3243), .Y(register__n8226) );
  BUFx4f_ASAP7_75t_R register___U4095 ( .A(register__n3244), .Y(register__n3243) );
  AND3x1_ASAP7_75t_R register___U4096 ( .A(register__n10590), .B(register__n10588), .C(register__n10589), .Y(register__n1281) );
  AND2x2_ASAP7_75t_R register___U4097 ( .A(register__n8693), .B(register__n1281), .Y(register__n7323) );
  INVxp33_ASAP7_75t_R register___U4098 ( .A(register__n572), .Y(register__n1282) );
  HB1xp67_ASAP7_75t_R register___U4099 ( .A(register__n12896), .Y(register__n3331) );
  AO22x1_ASAP7_75t_R register___U4100 ( .A1(register__net91021), .A2(register__net126316), .B1(register__net89741), 
        .B2(register__net123880), .Y(register__n11005) );
  AO22x1_ASAP7_75t_R register___U4101 ( .A1(register__n9617), .A2(register__net126316), .B1(register__n8947), .B2(
        net123880), .Y(register__n10580) );
  AO22x1_ASAP7_75t_R register___U4102 ( .A1(register__n9343), .A2(register__net126316), .B1(register__n9369), .B2(
        net123880), .Y(register__n11070) );
  AO22x1_ASAP7_75t_R register___U4103 ( .A1(register__n9611), .A2(register__net126316), .B1(register__n10078), .B2(
        net123880), .Y(register__n10921) );
  AO22x1_ASAP7_75t_R register___U4104 ( .A1(register__n9609), .A2(register__net126316), .B1(register__n10074), .B2(
        net123880), .Y(register__n10942) );
  AO22x1_ASAP7_75t_R register___U4105 ( .A1(register__n9812), .A2(register__net126316), .B1(register__n10142), .B2(
        net123880), .Y(register__n10747) );
  AO22x1_ASAP7_75t_R register___U4106 ( .A1(register__net90649), .A2(register__net126316), .B1(register__net100994), 
        .B2(register__net123880), .Y(register__n10708) );
  AO22x1_ASAP7_75t_R register___U4107 ( .A1(register__n9619), .A2(register__net126316), .B1(register__n10066), .B2(
        net123880), .Y(register__n10539) );
  AO22x1_ASAP7_75t_R register___U4108 ( .A1(register__n9853), .A2(register__net126316), .B1(register__n10301), .B2(
        net123880), .Y(register__n11026) );
  BUFx3_ASAP7_75t_R register___U4109 ( .A(register__n7651), .Y(register__n3184) );
  INVxp67_ASAP7_75t_R register___U4110 ( .A(register__n3764), .Y(register__n6175) );
  HB1xp67_ASAP7_75t_R register___U4111 ( .A(register__n3892), .Y(register__n3891) );
  XNOR2x2_ASAP7_75t_R register___U4112 ( .A(register__n1422), .B(register__n154), .Y(register__n12514) );
  AO22x1_ASAP7_75t_R register___U4113 ( .A1(register__n7988), .A2(register__net125170), .B1(register__n8799), .B2(register__n515), 
        .Y(register__n11529) );
  BUFx6f_ASAP7_75t_R register___U4114 ( .A(register__net112763), .Y(register__net66306) );
  AO22x1_ASAP7_75t_R register___U4115 ( .A1(register__n9692), .A2(register__C6423_net61340), .B1(register__n9963), .B2(
        net125365), .Y(register__n11233) );
  AO22x1_ASAP7_75t_R register___U4116 ( .A1(register__n9690), .A2(register__C6423_net61340), .B1(register__n9961), .B2(
        net125365), .Y(register__n11253) );
  AO22x1_ASAP7_75t_R register___U4117 ( .A1(register__n9694), .A2(register__C6423_net61340), .B1(register__n9965), .B2(
        net125365), .Y(register__n11212) );
  AO22x1_ASAP7_75t_R register___U4118 ( .A1(register__n7990), .A2(register__C6423_net61340), .B1(register__n9363), .B2(
        net125365), .Y(register__n11334) );
  AO22x1_ASAP7_75t_R register___U4119 ( .A1(register__n9768), .A2(register__C6423_net61340), .B1(register__n10110), 
        .B2(register__net125365), .Y(register__n11379) );
  AND2x4_ASAP7_75t_R register___U4120 ( .A(register__n11720), .B(register__n11728), .Y(register__net125365) );
  INVxp67_ASAP7_75t_R register___U4121 ( .A(register__n12580), .Y(register__n9394) );
  BUFx6f_ASAP7_75t_R register___U4122 ( .A(register__net115027), .Y(register__net115025) );
  BUFx12f_ASAP7_75t_R register___U4123 ( .A(register__n3877), .Y(register__n3839) );
  AO21x1_ASAP7_75t_R register___U4124 ( .A1(register__net91105), .A2(register__net117657), .B(register__n2400), .Y(
        n1285) );
  AO22x1_ASAP7_75t_R register___U4125 ( .A1(register__n12136), .A2(register__n1333), .B1(register__n1334), .B2(register__n1411), 
        .Y(register__n1286) );
  HB1xp67_ASAP7_75t_R register___U4126 ( .A(register__n12697), .Y(register__n4670) );
  AND3x1_ASAP7_75t_R register___U4127 ( .A(register__n11448), .B(register__n8751), .C(register__n11447), .Y(register__n1287) );
  AND2x2_ASAP7_75t_R register___U4128 ( .A(register__n7016), .B(register__n1287), .Y(register__n7887) );
  HB1xp67_ASAP7_75t_R register___U4129 ( .A(register__n12772), .Y(register__n3764) );
  AND2x2_ASAP7_75t_R register___U4130 ( .A(register__n2089), .B(register__n3240), .Y(register__n1290) );
  INVx2_ASAP7_75t_R register___U4131 ( .A(register__n3241), .Y(register__n6426) );
  AO22x1_ASAP7_75t_R register___U4132 ( .A1(register__n7810), .A2(register__net129746), .B1(register__n6877), .B2(
        net139537), .Y(register__n10795) );
  BUFx2_ASAP7_75t_R register___U4133 ( .A(register__n3242), .Y(register__n3241) );
  HB1xp67_ASAP7_75t_R register___U4134 ( .A(register__n13048), .Y(register__n3892) );
  INVxp67_ASAP7_75t_R register___U4135 ( .A(register__n10591), .Y(register__n8693) );
  INVxp67_ASAP7_75t_R register___U4136 ( .A(register__n13091), .Y(register__n4973) );
  INVxp33_ASAP7_75t_R register___U4137 ( .A(register__n4270), .Y(register__n1548) );
  HB1xp67_ASAP7_75t_R register___U4138 ( .A(register__n11634), .Y(register__n3242) );
  HB1xp67_ASAP7_75t_R register___U4139 ( .A(register__n3941), .Y(register__n2864) );
  AO22x1_ASAP7_75t_R register___U4140 ( .A1(register__n9284), .A2(register__n768), .B1(register__n10231), .B2(register__n75), .Y(
        n10752) );
  HB1xp67_ASAP7_75t_R register___U4141 ( .A(register__n11332), .Y(register__n5617) );
  HB1xp67_ASAP7_75t_R register___U4142 ( .A(register__n5617), .Y(register__n5616) );
  AO22x1_ASAP7_75t_R register___U4143 ( .A1(register__n8345), .A2(register__C6423_net61318), .B1(register__n10026), 
        .B2(register__n1448), .Y(register__n11250) );
  AO22x1_ASAP7_75t_R register___U4144 ( .A1(register__n8205), .A2(register__n128), .B1(register__n8550), .B2(register__n1454), 
        .Y(register__n11668) );
  AO22x1_ASAP7_75t_R register___U4145 ( .A1(register__n7680), .A2(register__C6423_net61318), .B1(register__n10201), 
        .B2(register__n1445), .Y(register__n11418) );
  AOI22xp33_ASAP7_75t_R register___U4146 ( .A1(register__n8797), .A2(register__net117658), .B1(register__n9132), .B2(
        n841), .Y(register__n1291) );
  AO22x1_ASAP7_75t_R register___U4147 ( .A1(register__n10477), .A2(register__net117657), .B1(register__n10456), .B2(
        n839), .Y(register__n10666) );
  BUFx4f_ASAP7_75t_R register___U4148 ( .A(register__n7701), .Y(register__n7700) );
  BUFx6f_ASAP7_75t_R register___U4149 ( .A(register__net66306), .Y(register__net66304) );
  INVx1_ASAP7_75t_R register___U4150 ( .A(register__n10997), .Y(register__n1292) );
  HB1xp67_ASAP7_75t_R register___U4151 ( .A(register__n12450), .Y(register__n6269) );
  AO22x1_ASAP7_75t_R register___U4152 ( .A1(register__net96895), .A2(register__net125170), .B1(register__net90077), 
        .B2(register__n235), .Y(register__n11267) );
  INVx1_ASAP7_75t_R register___U4153 ( .A(register__register__n12937), .Y(register__n1293) );
  AND2x2_ASAP7_75t_R register___U4154 ( .A(register__n10994), .B(register__n10996), .Y(register__n1294) );
  AND3x1_ASAP7_75t_R register___U4155 ( .A(register__n1294), .B(register__n10995), .C(register__n1292), .Y(register__n9178) );
  AOI22xp33_ASAP7_75t_R register___U4156 ( .A1(register__n4001), .A2(register__n1058), .B1(register__n1295), .B2(register__n103), 
        .Y(register__n13165) );
  CKINVDCx20_ASAP7_75t_R register___U4157 ( .A(register__n9567), .Y(register__n1295) );
  AOI22xp33_ASAP7_75t_R register___U4158 ( .A1(register__n4001), .A2(register__n3336), .B1(register__n1296), .B2(register__n1266), 
        .Y(register__n13135) );
  CKINVDCx20_ASAP7_75t_R register___U4159 ( .A(register__n9768), .Y(register__n1296) );
  OAI21xp33_ASAP7_75t_R register___U4160 ( .A1(register__n2592), .A2(register__n_cell_124679_net155985), .B(
        n2621), .Y(register__n2622) );
  BUFx4f_ASAP7_75t_R register___U4161 ( .A(register__n4966), .Y(register__n12238) );
  AO22x1_ASAP7_75t_R register___U4162 ( .A1(register__n6960), .A2(register__n39), .B1(register__n6624), .B2(
        C6422_net60399), .Y(register__n10687) );
  AO22x1_ASAP7_75t_R register___U4163 ( .A1(register__net104592), .A2(register__n39), .B1(register__net89409), .B2(
        C6422_net60399), .Y(register__n10808) );
  AO22x1_ASAP7_75t_R register___U4164 ( .A1(register__net91045), .A2(register__n39), .B1(register__net89877), .B2(
        C6422_net60399), .Y(register__n10873) );
  AO22x1_ASAP7_75t_R register___U4165 ( .A1(register__n8343), .A2(register__n39), .B1(register__n10020), .B2(
        C6422_net60399), .Y(register__n10919) );
  AO22x1_ASAP7_75t_R register___U4166 ( .A1(register__net90217), .A2(register__n39), .B1(register__net93661), .B2(
        C6422_net60399), .Y(register__n11087) );
  AO22x1_ASAP7_75t_R register___U4167 ( .A1(register__n9597), .A2(register__n39), .B1(register__n10018), .B2(
        C6422_net60399), .Y(register__n10963) );
  AO22x1_ASAP7_75t_R register___U4168 ( .A1(register__n10479), .A2(register__n39), .B1(register__n10452), .B2(register__net137523), .Y(register__n10940) );
  AO22x1_ASAP7_75t_R register___U4169 ( .A1(register__n9256), .A2(register__n40), .B1(register__n10028), .B2(
        C6422_net60399), .Y(register__n10578) );
  AO22x1_ASAP7_75t_R register___U4170 ( .A1(register__n9834), .A2(register__n40), .B1(register__n6645), .B2(
        C6422_net60399), .Y(register__n10984) );
  AO22x1_ASAP7_75t_R register___U4171 ( .A1(register__n7514), .A2(register__n39), .B1(register__n6630), .B2(
        C6422_net60399), .Y(register__n10645) );
  AO22x1_ASAP7_75t_R register___U4172 ( .A1(register__net104579), .A2(register__n39), .B1(register__net101048), .B2(
        C6422_net60399), .Y(register__n10706) );
  AO22x1_ASAP7_75t_R register___U4173 ( .A1(register__net106940), .A2(register__n40), .B1(register__net89889), .B2(
        C6422_net60399), .Y(register__n11003) );
  AO22x1_ASAP7_75t_R register___U4174 ( .A1(register__n9840), .A2(register__n39), .B1(register__n8171), .B2(
        C6422_net60399), .Y(register__n11045) );
  AO22x1_ASAP7_75t_R register___U4175 ( .A1(register__n7992), .A2(register__n39), .B1(register__n10307), .B2(
        C6422_net60399), .Y(register__n10850) );
  AO22x1_ASAP7_75t_R register___U4176 ( .A1(register__n8345), .A2(register__n39), .B1(register__n10026), .B2(
        C6422_net60399), .Y(register__n10623) );
  AO22x1_ASAP7_75t_R register___U4177 ( .A1(register__n9601), .A2(register__n39), .B1(register__n10024), .B2(
        C6422_net60399), .Y(register__n10668) );
  AO22x1_ASAP7_75t_R register___U4178 ( .A1(register__n7680), .A2(register__n40), .B1(register__n10201), .B2(
        C6422_net60399), .Y(register__n10792) );
  AO22x1_ASAP7_75t_R register___U4179 ( .A1(register__n8206), .A2(register__n39), .B1(register__n8549), .B2(
        C6422_net60399), .Y(register__n11068) );
  HB1xp67_ASAP7_75t_R register___U4180 ( .A(register__n11944), .Y(register__n11938) );
  BUFx2_ASAP7_75t_R register___U4181 ( .A(register__n10839), .Y(register__n5915) );
  AND4x2_ASAP7_75t_R register___U4182 ( .A(register__n4760), .B(register__n33), .C(register__n4761), .D(register__n3060), .Y(
        n10840) );
  INVx1_ASAP7_75t_R register___U4183 ( .A(register__n10629), .Y(register__n1298) );
  NAND3xp33_ASAP7_75t_R register___U4184 ( .A(register__n1954), .B(register__n429), .C(IF_ID_rs1[2]), 
        .Y(register__n1299) );
  INVx1_ASAP7_75t_R register___U4185 ( .A(register__n11240), .Y(register__n1316) );
  HB1xp67_ASAP7_75t_R register___U4186 ( .A(register__n5027), .Y(register__n5026) );
  HB1xp67_ASAP7_75t_R register___U4187 ( .A(register__n11144), .Y(register__n5027) );
  INVxp67_ASAP7_75t_R register___U4188 ( .A(register__n2927), .Y(register__n4380) );
  HB1xp67_ASAP7_75t_R register___U4189 ( .A(register__n10791), .Y(register__n2927) );
  HB1xp67_ASAP7_75t_R register___U4190 ( .A(register__n5168), .Y(register__n5167) );
  HB1xp67_ASAP7_75t_R register___U4191 ( .A(register__n11014), .Y(register__n5168) );
  INVx1_ASAP7_75t_R register___U4192 ( .A(register__n10609), .Y(register__n1300) );
  NOR3x1_ASAP7_75t_R register___U4193 ( .A(register__n1484), .B(register__n4622), .C(register__n8257), .Y(register__n11680) );
  INVxp33_ASAP7_75t_R register___U4194 ( .A(register__n4335), .Y(register__n7322) );
  BUFx6f_ASAP7_75t_R register___U4195 ( .A(register__n7592), .Y(register__n8619) );
  INVxp67_ASAP7_75t_R register___U4196 ( .A(register__n4707), .Y(register__n7270) );
  BUFx12f_ASAP7_75t_R register___U4197 ( .A(register__net112764), .Y(register__net112762) );
  AO22x1_ASAP7_75t_R register___U4198 ( .A1(register__n6850), .A2(register__n38), .B1(register__n10460), .B2(register__n366), .Y(
        n10565) );
  AOI21xp33_ASAP7_75t_R register___U4199 ( .A1(register__net123879), .A2(register__net89717), .B(register__n2388), .Y(
        n2407) );
  OA22x2_ASAP7_75t_R register___U4200 ( .A1(register__net64414), .A2(register__n1301), .B1(register__net88496), .B2(
        n1302), .Y(register__n12908) );
  HB1xp67_ASAP7_75t_R register___U4201 ( .A(register__n12808), .Y(register__n3588) );
  INVxp67_ASAP7_75t_R register___U4202 ( .A(register__n3046), .Y(register__n4770) );
  HB1xp67_ASAP7_75t_R register___U4203 ( .A(register__n3047), .Y(register__n3046) );
  AOI21xp33_ASAP7_75t_R register___U4204 ( .A1(register__net120788), .A2(register__net90961), .B(register__n2365), .Y(
        n2367) );
  AO22x1_ASAP7_75t_R register___U4205 ( .A1(register__n9863), .A2(register__net120788), .B1(register__n7230), .B2(register__n369), 
        .Y(register__n10693) );
  AO22x1_ASAP7_75t_R register___U4206 ( .A1(register__net96863), .A2(register__C6422_net60445), .B1(register__net107943), .B2(register__C6422_net60443), .Y(register__n10712) );
  AO22x1_ASAP7_75t_R register___U4207 ( .A1(register__n9627), .A2(register__n38), .B1(register__n10090), .B2(
        C6422_net60443), .Y(register__n10674) );
  CKINVDCx20_ASAP7_75t_R register___U4208 ( .A(register__n9836), .Y(register__n1307) );
  CKINVDCx20_ASAP7_75t_R register___U4209 ( .A(register__n5929), .Y(register__n1308) );
  AO22x1_ASAP7_75t_R register___U4210 ( .A1(register__n9095), .A2(register__net110414), .B1(register__n10165), .B2(
        net117889), .Y(register__n11634) );
  INVx2_ASAP7_75t_R register___U4211 ( .A(register__net112762), .Y(register__n1467) );
  HB1xp67_ASAP7_75t_R register___U4212 ( .A(register__n12506), .Y(register__n7679) );
  AO22x1_ASAP7_75t_R register___U4213 ( .A1(register__net64456), .A2(register__n2020), .B1(register__n1311), .B2(register__n1312), 
        .Y(register__n1310) );
  CKINVDCx20_ASAP7_75t_R register___U4214 ( .A(register__net100992), .Y(register__n1311) );
  CKINVDCx14_ASAP7_75t_R register___U4215 ( .A(register__n2020), .Y(register__n1989) );
  NOR2xp33_ASAP7_75t_R register___U4216 ( .A(register__n11602), .B(register__n1324), .Y(register__n1387) );
  INVx1_ASAP7_75t_R register___U4217 ( .A(register__n10636), .Y(register__n1315) );
  NOR4xp75_ASAP7_75t_R register___U4218 ( .A(register__n1316), .B(register__n5995), .C(register__n1317), .D(register__n1318), .Y(
        n9155) );
  NAND4xp75_ASAP7_75t_R register___U4219 ( .A(register__n7307), .B(register__n1516), .C(register__n6750), .D(register__n4609), 
        .Y(register__n1317) );
  INVx6_ASAP7_75t_R register___U4220 ( .A(register__n12303), .Y(register__n12288) );
  BUFx12f_ASAP7_75t_R register___U4221 ( .A(register__n4815), .Y(register__n12303) );
  INVx1_ASAP7_75t_R register___U4222 ( .A(register__n10841), .Y(register__n7976) );
  AO22x1_ASAP7_75t_R register___U4223 ( .A1(register__n9881), .A2(register__net110414), .B1(register__n10321), .B2(
        n1129), .Y(register__n11468) );
  HB1xp67_ASAP7_75t_R register___U4224 ( .A(register__n11509), .Y(register__n4707) );
  HB1xp67_ASAP7_75t_R register___U4225 ( .A(register__net63390), .Y(register__net63358) );
  HB1xp67_ASAP7_75t_R register___U4226 ( .A(register__net63390), .Y(register__net63354) );
  HB1xp67_ASAP7_75t_R register___U4227 ( .A(register__net63390), .Y(register__net63360) );
  HB1xp67_ASAP7_75t_R register___U4228 ( .A(register__net63390), .Y(register__net63356) );
  INVx1_ASAP7_75t_R register___U4229 ( .A(register__net63358), .Y(register__net63326) );
  INVx1_ASAP7_75t_R register___U4230 ( .A(register__net63354), .Y(register__net63320) );
  INVx1_ASAP7_75t_R register___U4231 ( .A(register__net63360), .Y(register__net63328) );
  INVx1_ASAP7_75t_R register___U4232 ( .A(register__net63356), .Y(register__net63322) );
  INVxp67_ASAP7_75t_R register___U4233 ( .A(register__net64784), .Y(register__net64750) );
  HB1xp67_ASAP7_75t_R register___U4234 ( .A(register__n2837), .Y(register__n2836) );
  INVxp67_ASAP7_75t_R register___U4235 ( .A(register__n2836), .Y(register__n3869) );
  INVxp67_ASAP7_75t_R register___U4236 ( .A(register__n12579), .Y(register__n5372) );
  INVxp33_ASAP7_75t_R register___U4237 ( .A(register__n4270), .Y(register__n2078) );
  HB1xp67_ASAP7_75t_R register___U4238 ( .A(register__net64818), .Y(register__net64804) );
  HB1xp67_ASAP7_75t_R register___U4239 ( .A(register__net64818), .Y(register__net64802) );
  BUFx6f_ASAP7_75t_R register___U4240 ( .A(register__net64788), .Y(register__net144464) );
  INVx1_ASAP7_75t_R register___U4241 ( .A(register__n11377), .Y(register__n1319) );
  BUFx6f_ASAP7_75t_R register___U4242 ( .A(register__net130079), .Y(register__net95787) );
  BUFx6f_ASAP7_75t_R register___U4243 ( .A(register__net95787), .Y(register__C6423_net69178) );
  OA22x2_ASAP7_75t_R register___U4244 ( .A1(register__net64424), .A2(register__n460), .B1(register__n1320), .B2(register__n472), 
        .Y(register__n12939) );
  CKINVDCx20_ASAP7_75t_R register___U4245 ( .A(register__n1763), .Y(register__n1320) );
  INVx6_ASAP7_75t_R register___U4246 ( .A(register__net64456), .Y(register__net64424) );
  HB1xp67_ASAP7_75t_R register___U4247 ( .A(register__net123601), .Y(register__net64806) );
  AO22x1_ASAP7_75t_R register___U4248 ( .A1(register__n8160), .A2(register__C6423_net61343), .B1(register__n10158), 
        .B2(register__net129787), .Y(register__n11509) );
  AO22x1_ASAP7_75t_R register___U4249 ( .A1(register__n9628), .A2(register__n38), .B1(register__n10091), .B2(register__n369), .Y(
        n10629) );
  AO22x1_ASAP7_75t_R register___U4250 ( .A1(register__n9903), .A2(register__net138040), .B1(register__n10206), .B2(
        net125803), .Y(register__n11691) );
  AO22x1_ASAP7_75t_R register___U4251 ( .A1(register__n9664), .A2(register__net125426), .B1(register__n9993), .B2(
        net125804), .Y(register__n11251) );
  INVx1_ASAP7_75t_R register___U4252 ( .A(register__net138525), .Y(register__net64754) );
  HB1xp67_ASAP7_75t_R register___U4253 ( .A(register__net64804), .Y(register__net138525) );
  INVx1_ASAP7_75t_R register___U4254 ( .A(register__n11424), .Y(register__n7598) );
  AO22x1_ASAP7_75t_R register___U4255 ( .A1(register__n9853), .A2(register__C6423_net61343), .B1(register__n10301), 
        .B2(register__net129787), .Y(register__n11630) );
  AO22x1_ASAP7_75t_R register___U4256 ( .A1(register__n9911), .A2(register__n413), .B1(register__n10214), .B2(register__net126602), .Y(register__n10791) );
  HB1xp67_ASAP7_75t_R register___U4257 ( .A(register__n12309), .Y(register__n4746) );
  BUFx2_ASAP7_75t_R register___U4258 ( .A(register__n4717), .Y(register__n4716) );
  BUFx12f_ASAP7_75t_R register___U4259 ( .A(register__net91919), .Y(register__net142364) );
  INVx1_ASAP7_75t_R register___U4260 ( .A(register__n11274), .Y(register__n1323) );
  NAND4xp25_ASAP7_75t_R register___U4261 ( .A(register__n4729), .B(register__n7066), .C(register__n6412), .D(register__n7065), 
        .Y(register__n1324) );
  INVx1_ASAP7_75t_R register___U4262 ( .A(register__n11333), .Y(register__n1325) );
  AO22x1_ASAP7_75t_R register___U4263 ( .A1(register__n6849), .A2(register__net110414), .B1(register__n10460), .B2(
        n1074), .Y(register__n11192) );
  AO22x1_ASAP7_75t_R register___U4264 ( .A1(register__n9634), .A2(register__C6423_net69526), .B1(register__n7477), .B2(
        n1074), .Y(register__n11170) );
  INVxp67_ASAP7_75t_R register___U4265 ( .A(register__n12554), .Y(register__n7025) );
  BUFx6f_ASAP7_75t_R register___U4266 ( .A(register__n3374), .Y(register__n1326) );
  AO22x1_ASAP7_75t_R register___U4267 ( .A1(register__n9734), .A2(register__C6422_net60408), .B1(register__n8511), .B2(
        n835), .Y(register__n10982) );
  OAI22xp5_ASAP7_75t_R register___U4268 ( .A1(register__n53), .A2(register__n8642), .B1(register__net61369), .B2(register__n12466), .Y(read_reg_data_1[30]) );
  AO22x1_ASAP7_75t_R register___U4269 ( .A1(register__n7193), .A2(register__C6423_net61343), .B1(register__n10273), 
        .B2(register__net129787), .Y(register__n11358) );
  AO22x1_ASAP7_75t_R register___U4270 ( .A1(register__n9343), .A2(register__C6423_net61343), .B1(register__n9369), .B2(
        net122313), .Y(register__n11670) );
  INVx2_ASAP7_75t_R register___U4271 ( .A(register__n7700), .Y(register__n9191) );
  BUFx3_ASAP7_75t_R register___U4272 ( .A(register__n11101), .Y(register__n7701) );
  INVx1_ASAP7_75t_R register___U4273 ( .A(register__n11269), .Y(register__n1328) );
  HB1xp67_ASAP7_75t_R register___U4274 ( .A(register__n1291), .Y(register__n3063) );
  INVxp67_ASAP7_75t_R register___U4275 ( .A(register__n10637), .Y(register__n8310) );
  AND2x2_ASAP7_75t_R register___U4276 ( .A(register__n8013), .B(register__n1502), .Y(register__n1329) );
  NAND4xp25_ASAP7_75t_R register___U4277 ( .A(register__n20), .B(register__n4483), .C(register__n4978), .D(register__n1648), .Y(
        n1330) );
  BUFx6f_ASAP7_75t_R register___U4278 ( .A(register__n3004), .Y(register__n3069) );
  HB1xp67_ASAP7_75t_R register___U4279 ( .A(register__n12416), .Y(register__n3569) );
  BUFx12f_ASAP7_75t_R register___U4280 ( .A(register__n1997), .Y(register__net130666) );
  NAND4xp25_ASAP7_75t_R register___U4281 ( .A(register__n8270), .B(register__n8269), .C(register__n9170), .D(register__n8268), 
        .Y(register__n2245) );
  INVx1_ASAP7_75t_R register___U4282 ( .A(register__n11591), .Y(register__n8268) );
  OAI22xp33_ASAP7_75t_R register___U4283 ( .A1(register__n1331), .A2(register__C6423_net72243), .B1(register__n1332), 
        .B2(register__n_cell_124679_net155985), .Y(register__n11210) );
  CKINVDCx20_ASAP7_75t_R register___U4284 ( .A(register__n9666), .Y(register__n1331) );
  CKINVDCx20_ASAP7_75t_R register___U4285 ( .A(register__n9425), .Y(register__n1332) );
  INVx4_ASAP7_75t_R register___U4286 ( .A(register__n12253), .Y(register__n1910) );
  INVx6_ASAP7_75t_R register___U4287 ( .A(register__n12267), .Y(register__n12253) );
  AOI211x1_ASAP7_75t_R register___U4288 ( .A1(register__net126316), .A2(register__net90261), .B(register__n2677), .C(
        n2653), .Y(register__n2676) );
  CKINVDCx20_ASAP7_75t_R register___U4289 ( .A(register__n8753), .Y(register__n1334) );
  INVx4_ASAP7_75t_R register___U4290 ( .A(register__n1411), .Y(register__n1419) );
  HB1xp67_ASAP7_75t_R register___U4291 ( .A(register__n13000), .Y(register__n5271) );
  INVxp67_ASAP7_75t_R register___U4292 ( .A(register__n5272), .Y(register__n6190) );
  INVxp33_ASAP7_75t_R register___U4293 ( .A(register__n4682), .Y(register__n7925) );
  INVxp67_ASAP7_75t_R register___U4294 ( .A(register__n12135), .Y(register__n12119) );
  HB1xp67_ASAP7_75t_R register___U4295 ( .A(register__n7925), .Y(register__n4683) );
  HB1xp67_ASAP7_75t_R register___U4296 ( .A(register__n11948), .Y(register__n11941) );
  HB1xp67_ASAP7_75t_R register___U4297 ( .A(register__n11948), .Y(register__n11942) );
  AO22x1_ASAP7_75t_R register___U4298 ( .A1(register__n10483), .A2(register__C6423_net61343), .B1(register__n10463), 
        .B2(register__net122313), .Y(register__n11333) );
  HB1xp67_ASAP7_75t_R register___U4299 ( .A(register__n8607), .Y(register__n6803) );
  INVxp67_ASAP7_75t_R register___U4300 ( .A(register__n3783), .Y(register__n5383) );
  INVx6_ASAP7_75t_R register___U4301 ( .A(register__n12131), .Y(register__n12116) );
  BUFx12f_ASAP7_75t_R register___U4302 ( .A(register__n12135), .Y(register__n12131) );
  INVxp67_ASAP7_75t_R register___U4303 ( .A(register__n5101), .Y(register__n5911) );
  NOR4xp75_ASAP7_75t_R register___U4304 ( .A(register__n3228), .B(register__n3229), .C(register__n11339), .D(register__n11340), 
        .Y(register__n11320) );
  BUFx3_ASAP7_75t_R register___U4305 ( .A(register__n11337), .Y(register__n3228) );
  BUFx3_ASAP7_75t_R register___U4306 ( .A(register__n11338), .Y(register__n3229) );
  AO22x1_ASAP7_75t_R register___U4307 ( .A1(register__n9648), .A2(register__net109849), .B1(register__n9975), .B2(register__n632), 
        .Y(register__n11340) );
  HB1xp67_ASAP7_75t_R register___U4308 ( .A(register__n11982), .Y(register__n3020) );
  HB1xp67_ASAP7_75t_R register___U4309 ( .A(register__n3784), .Y(register__n3783) );
  BUFx6f_ASAP7_75t_R register___U4310 ( .A(register__n5348), .Y(register__n5344) );
  INVxp67_ASAP7_75t_R register___U4311 ( .A(register__n13158), .Y(register__n6434) );
  NOR2xp33_ASAP7_75t_R register___U4312 ( .A(register__n368), .B(register__n1338), .Y(register__n1339) );
  NOR2xp33_ASAP7_75t_R register___U4313 ( .A(register__n1339), .B(register__n2363), .Y(register__n2320) );
  INVxp33_ASAP7_75t_R register___U4314 ( .A(register__net89685), .Y(register__n1338) );
  BUFx6f_ASAP7_75t_R register___U4315 ( .A(register__net89686), .Y(register__net89685) );
  INVxp33_ASAP7_75t_R register___U4316 ( .A(register__n5548), .Y(register__n1646) );
  INVxp33_ASAP7_75t_R register___U4317 ( .A(register__n5548), .Y(register__n1645) );
  INVxp33_ASAP7_75t_R register___U4318 ( .A(register__n5548), .Y(register__n1644) );
  INVx1_ASAP7_75t_R register___U4319 ( .A(register__n11231), .Y(register__n1340) );
  AO22x1_ASAP7_75t_R register___U4320 ( .A1(register__n7801), .A2(register__net93569), .B1(register__n8134), .B2(
        net147379), .Y(register__n11318) );
  HB1xp67_ASAP7_75t_R register___U4321 ( .A(register__n11210), .Y(register__n4682) );
  NOR4xp25_ASAP7_75t_R register___U4322 ( .A(register__n11677), .B(register__n3211), .C(register__n2878), .D(register__n11674), 
        .Y(register__n11657) );
  AO22x1_ASAP7_75t_R register___U4323 ( .A1(register__n10505), .A2(register__n481), .B1(register__n10425), .B2(register__n633), 
        .Y(register__n11677) );
  BUFx3_ASAP7_75t_R register___U4324 ( .A(register__n11675), .Y(register__n3211) );
  BUFx3_ASAP7_75t_R register___U4325 ( .A(register__n11676), .Y(register__n2878) );
  HB1xp67_ASAP7_75t_R register___U4326 ( .A(register__n4336), .Y(register__n4335) );
  INVx1_ASAP7_75t_R register___U4327 ( .A(register__n11576), .Y(register__n1341) );
  NAND2xp33_ASAP7_75t_R register___U4328 ( .A(register__n1342), .B(register__n1851), .Y(register__n1343) );
  INVxp33_ASAP7_75t_R register___U4329 ( .A(register__net63276), .Y(register__n1342) );
  INVxp67_ASAP7_75t_R register___U4330 ( .A(register__n4144), .Y(register__n5219) );
  AO22x1_ASAP7_75t_R register___U4331 ( .A1(register__net90961), .A2(register__net110414), .B1(register__net89685), 
        .B2(register__n1073), .Y(register__n11274) );
  INVx1_ASAP7_75t_R register___U4332 ( .A(register__n1345), .Y(register__n1350) );
  AOI21xp33_ASAP7_75t_R register___U4333 ( .A1(register__n387), .A2(register__net90733), .B(register__n2383), .Y(register__n2403)
         );
  AO22x1_ASAP7_75t_R register___U4334 ( .A1(register__n9897), .A2(register__net131160), .B1(register__n10223), .B2(
        net120912), .Y(register__n11072) );
  AO22x1_ASAP7_75t_R register___U4335 ( .A1(register__net90457), .A2(register__net131160), .B1(register__net89209), 
        .B2(register__net120912), .Y(register__n10710) );
  AO22x1_ASAP7_75t_R register___U4336 ( .A1(register__n7704), .A2(register__net131160), .B1(register__n8030), .B2(
        net120912), .Y(register__n10967) );
  AO22x1_ASAP7_75t_R register___U4337 ( .A1(register__n8911), .A2(register__net131160), .B1(register__n10048), .B2(
        net120912), .Y(register__n10582) );
  AO22x1_ASAP7_75t_R register___U4338 ( .A1(register__n9732), .A2(register__n387), .B1(register__n10303), .B2(register__n326), 
        .Y(register__n11028) );
  BUFx12f_ASAP7_75t_R register___U4339 ( .A(register__n3668), .Y(register__n7610) );
  AO22x1_ASAP7_75t_R register___U4340 ( .A1(register__n9804), .A2(register__net93569), .B1(register__n10203), .B2(register__n284), 
        .Y(register__n11698) );
  AO22x1_ASAP7_75t_R register___U4341 ( .A1(register__n9830), .A2(register__net110414), .B1(register__n10271), .B2(
        n1074), .Y(register__n11596) );
  HB1xp67_ASAP7_75t_R register___U4342 ( .A(register__n11724), .Y(register__n3078) );
  AO22x1_ASAP7_75t_R register___U4343 ( .A1(register__n9861), .A2(register__n309), .B1(register__n10295), .B2(register__net147378), .Y(register__n11724) );
  HB1xp67_ASAP7_75t_R register___U4344 ( .A(register__n5102), .Y(register__n5101) );
  HB1xp67_ASAP7_75t_R register___U4345 ( .A(WB_rd[1]), .Y(register__n5523) );
  INVxp33_ASAP7_75t_R register___U4346 ( .A(register__n3093), .Y(register__n7012) );
  INVxp67_ASAP7_75t_R register___U4347 ( .A(register__n6493), .Y(register__n6826) );
  OAI22xp5_ASAP7_75t_R register___U4348 ( .A1(register__n53), .A2(register__n4032), .B1(register__net61369), .B2(register__n12264), .Y(read_reg_data_1[18]) );
  INVxp67_ASAP7_75t_R register___U4349 ( .A(register__n3127), .Y(register__n6197) );
  HB1xp67_ASAP7_75t_R register___U4350 ( .A(register__n3128), .Y(register__n3127) );
  INVx2_ASAP7_75t_R register___U4351 ( .A(register__n7314), .Y(register__n1478) );
  INVx2_ASAP7_75t_R register___U4352 ( .A(register__n5619), .Y(register__n7314) );
  HB1xp67_ASAP7_75t_R register___U4353 ( .A(register__n5043), .Y(register__n12185) );
  HB1xp67_ASAP7_75t_R register___U4354 ( .A(register__n7012), .Y(register__n3094) );
  HB1xp67_ASAP7_75t_R register___U4355 ( .A(register__n10601), .Y(register__n3128) );
  AO22x1_ASAP7_75t_R register___U4356 ( .A1(register__n6839), .A2(register__net126316), .B1(register__n10072), .B2(
        net123880), .Y(register__n10965) );
  AO22x1_ASAP7_75t_R register___U4357 ( .A1(register__n7521), .A2(register__net93282), .B1(register__n10136), .B2(
        net125803), .Y(register__n11669) );
  NAND2xp67_ASAP7_75t_R register___U4358 ( .A(register__n1955), .B(register__n1956), .Y(register__n2740) );
  INVx2_ASAP7_75t_R register___U4359 ( .A(register__n7350), .Y(register__n8279) );
  INVx1_ASAP7_75t_R register___U4360 ( .A(register__n12924), .Y(register__n1362) );
  HB1xp67_ASAP7_75t_R register___U4361 ( .A(register__n6494), .Y(register__n6493) );
  AO22x1_ASAP7_75t_R register___U4362 ( .A1(register__n12478), .A2(register__n690), .B1(register__n1364), .B2(register__n702), 
        .Y(register__n1363) );
  CKINVDCx20_ASAP7_75t_R register___U4363 ( .A(register__n9555), .Y(register__n1364) );
  INVxp33_ASAP7_75t_R register___U4364 ( .A(register__n4851), .Y(register__n1843) );
  NAND2xp5_ASAP7_75t_R register___U4365 ( .A(register__n49), .B(register__n2160), .Y(register__n1365) );
  NAND2x1p5_ASAP7_75t_R register___U4366 ( .A(register__n1851), .B(register__n11990), .Y(register__n1366) );
  INVx1_ASAP7_75t_R register___U4367 ( .A(register__n12006), .Y(register__n11990) );
  NOR4xp25_ASAP7_75t_R register___U4368 ( .A(register__n10561), .B(register__n10562), .C(register__n10563), .D(register__n10564), 
        .Y(register__n10548) );
  BUFx6f_ASAP7_75t_R register___U4369 ( .A(register__net145200), .Y(register__net144161) );
  BUFx3_ASAP7_75t_R register___U4370 ( .A(register__n3170), .Y(register__n3391) );
  INVxp67_ASAP7_75t_R register___U4371 ( .A(register__n1718), .Y(register__n1719) );
  INVxp67_ASAP7_75t_R register___U4372 ( .A(register__n1720), .Y(register__n1721) );
  OAI22xp33_ASAP7_75t_R register___U4373 ( .A1(register__net64854), .A2(register__n337), .B1(register__net90961), .B2(
        n344), .Y(register__n1367) );
  HB1xp67_ASAP7_75t_R register___U4374 ( .A(register__net64864), .Y(register__net64878) );
  BUFx3_ASAP7_75t_R register___U4375 ( .A(register__n10572), .Y(register__n7360) );
  INVx2_ASAP7_75t_R register___U4376 ( .A(register__n7359), .Y(register__n9188) );
  INVx6_ASAP7_75t_R register___U4377 ( .A(register__n12098), .Y(register__n12086) );
  AOI22xp33_ASAP7_75t_R register___U4378 ( .A1(register__n8539), .A2(register__n1867), .B1(register__n7562), .B2(register__n1347), 
        .Y(register__n1368) );
  OAI21xp33_ASAP7_75t_R register___U4379 ( .A1(register__n2684), .A2(register__n2685), .B(register__n50), .Y(register__n2634) );
  INVxp67_ASAP7_75t_R register___U4380 ( .A(register__n1878), .Y(register__n13312) );
  HB1xp67_ASAP7_75t_R register___U4381 ( .A(register__n12762), .Y(register__n3903) );
  INVx2_ASAP7_75t_R register___U4382 ( .A(register__n3456), .Y(register__n1788) );
  HB1xp67_ASAP7_75t_R register___U4383 ( .A(register__net64878), .Y(register__net64868) );
  INVxp67_ASAP7_75t_R register___U4384 ( .A(register__n3460), .Y(register__n4769) );
  HB1xp67_ASAP7_75t_R register___U4385 ( .A(register__n3461), .Y(register__n3460) );
  CKINVDCx10_ASAP7_75t_R register___U4386 ( .A(register__n11873), .Y(register__n5515) );
  INVx2_ASAP7_75t_R register___U4387 ( .A(register__n10977), .Y(register__n7677) );
  HB1xp67_ASAP7_75t_R register___U4388 ( .A(register__n1368), .Y(register__n3060) );
  BUFx6f_ASAP7_75t_R register___U4389 ( .A(register__net143365), .Y(register__net64870) );
  CKINVDCx10_ASAP7_75t_R register___U4390 ( .A(register__net63166), .Y(register__net132155) );
  HB1xp67_ASAP7_75t_R register___U4391 ( .A(register__n10923), .Y(register__n6494) );
  AO22x1_ASAP7_75t_R register___U4392 ( .A1(register__n9706), .A2(register__n387), .B1(register__n10036), .B2(register__net120912), .Y(register__n10923) );
  HB1xp67_ASAP7_75t_R register___U4393 ( .A(register__n13324), .Y(register__n4522) );
  INVx1_ASAP7_75t_R register___U4394 ( .A(register__n11439), .Y(register__n1369) );
  AND2x2_ASAP7_75t_R register___U4395 ( .A(register__n8271), .B(register__n479), .Y(register__n1370) );
  INVx2_ASAP7_75t_R register___U4396 ( .A(register__n4021), .Y(register__n1433) );
  AO22x1_ASAP7_75t_R register___U4397 ( .A1(register__n9329), .A2(register__net117657), .B1(register__n7468), .B2(register__n834), 
        .Y(register__n10557) );
  AO22x1_ASAP7_75t_R register___U4398 ( .A1(register__n9577), .A2(register__C6422_net60408), .B1(register__n10062), 
        .B2(register__n835), .Y(register__n10535) );
  HB1xp67_ASAP7_75t_R register___U4399 ( .A(register__net124440), .Y(register__net124439) );
  HB1xp67_ASAP7_75t_R register___U4400 ( .A(register__net64878), .Y(register__net143365) );
  OAI22xp33_ASAP7_75t_R register___U4401 ( .A1(register__n1371), .A2(register__n1398), .B1(register__n1372), .B2(register__n833), 
        .Y(register__n10622) );
  CKINVDCx20_ASAP7_75t_R register___U4402 ( .A(register__n9254), .Y(register__n1371) );
  CKINVDCx20_ASAP7_75t_R register___U4403 ( .A(register__n10058), .Y(register__n1372) );
  HB1xp67_ASAP7_75t_R register___U4404 ( .A(register__n12584), .Y(register__n3429) );
  INVxp33_ASAP7_75t_R register___U4405 ( .A(register__n7633), .Y(register__n1808) );
  INVxp33_ASAP7_75t_R register___U4406 ( .A(register__n7633), .Y(register__n1810) );
  INVxp33_ASAP7_75t_R register___U4407 ( .A(register__n7633), .Y(register__n1809) );
  INVxp67_ASAP7_75t_R register___U4408 ( .A(register__n6236), .Y(register__n7283) );
  HB1xp67_ASAP7_75t_R register___U4409 ( .A(register__n6237), .Y(register__n6236) );
  INVxp67_ASAP7_75t_R register___U4410 ( .A(register__n4781), .Y(register__n5907) );
  HB1xp67_ASAP7_75t_R register___U4411 ( .A(register__n4782), .Y(register__n4781) );
  OAI21x1_ASAP7_75t_R register___U4412 ( .A1(register__net127380), .A2(register__n2376), .B(register__n1900), .Y(register__n2399)
         );
  INVxp67_ASAP7_75t_R register___U4413 ( .A(register__n12771), .Y(register__n6174) );
  BUFx2_ASAP7_75t_R register___U4414 ( .A(register__n4577), .Y(register__n12273) );
  NAND2xp33_ASAP7_75t_R register___U4415 ( .A(register__n5213), .B(register__n1105), .Y(register__n1377) );
  NAND2xp33_ASAP7_75t_R register___U4416 ( .A(register__n1377), .B(register__n1378), .Y(register__n11426) );
  HB1xp67_ASAP7_75t_R register___U4417 ( .A(register__n9806), .Y(register__n5213) );
  BUFx12f_ASAP7_75t_R register___U4418 ( .A(register__n7811), .Y(register__n10205) );
  HB1xp67_ASAP7_75t_R register___U4419 ( .A(register__n285), .Y(register__net147379) );
  AO22x1_ASAP7_75t_R register___U4420 ( .A1(register__n9704), .A2(register__n387), .B1(register__n10034), .B2(register__net120912), .Y(register__n10944) );
  AO22x1_ASAP7_75t_R register___U4421 ( .A1(register__net94803), .A2(register__n387), .B1(register__net89445), .B2(
        net120912), .Y(register__n11091) );
  AO22x1_ASAP7_75t_R register___U4422 ( .A1(register__n9700), .A2(register__n387), .B1(register__n10050), .B2(register__net120912), .Y(register__n10541) );
  AO22x1_ASAP7_75t_R register___U4423 ( .A1(register__n10499), .A2(register__n387), .B1(register__n10454), .B2(
        net120912), .Y(register__n10563) );
  HB1xp67_ASAP7_75t_R register___U4424 ( .A(register__n12882), .Y(register__n3431) );
  CKINVDCx20_ASAP7_75t_R register___U4425 ( .A(register__n10122), .Y(register__n1380) );
  INVxp33_ASAP7_75t_R register___U4426 ( .A(register__n2871), .Y(register__n3722) );
  INVxp67_ASAP7_75t_R register___U4427 ( .A(register__n13200), .Y(register__n6126) );
  BUFx6f_ASAP7_75t_R register___U4428 ( .A(register__n12065), .Y(register__n12072) );
  INVx1_ASAP7_75t_R register___U4429 ( .A(register__n12069), .Y(register__n12056) );
  AO22x1_ASAP7_75t_R register___U4430 ( .A1(register__n8755), .A2(register__C6422_net60408), .B1(register__n10060), 
        .B2(register__n838), .Y(register__n10601) );
  AO22x1_ASAP7_75t_R register___U4431 ( .A1(register__n9575), .A2(register__C6422_net60408), .B1(register__n9431), .B2(
        n839), .Y(register__n10576) );
  HB1xp67_ASAP7_75t_R register___U4432 ( .A(register__n5770), .Y(register__n4002) );
  HB1xp67_ASAP7_75t_R register___U4433 ( .A(register__net63384), .Y(register__net63382) );
  INVxp67_ASAP7_75t_R register___U4434 ( .A(register__n4425), .Y(register__n5947) );
  HB1xp67_ASAP7_75t_R register___U4435 ( .A(register__n4426), .Y(register__n4425) );
  INVxp67_ASAP7_75t_R register___U4436 ( .A(register__n3164), .Y(register__n7049) );
  HB1xp67_ASAP7_75t_R register___U4437 ( .A(register__n3165), .Y(register__n3164) );
  INVxp67_ASAP7_75t_R register___U4438 ( .A(register__n4918), .Y(register__n7069) );
  INVx1_ASAP7_75t_R register___U4439 ( .A(register__n12826), .Y(register__n1383) );
  HB1xp67_ASAP7_75t_R register___U4440 ( .A(register__n12795), .Y(register__n6237) );
  HB1xp67_ASAP7_75t_R register___U4441 ( .A(register__n3722), .Y(register__n2873) );
  HB1xp67_ASAP7_75t_R register___U4442 ( .A(register__net36441), .Y(register__net124440) );
  NOR2xp33_ASAP7_75t_R register___U4443 ( .A(register__n2309), .B(register__n1885), .Y(register__net36441) );
  HB1xp67_ASAP7_75t_R register___U4444 ( .A(register__n5273), .Y(register__n5272) );
  CKINVDCx20_ASAP7_75t_R register___U4445 ( .A(register__n9742), .Y(register__n1384) );
  INVx13_ASAP7_75t_R register___U4446 ( .A(register__n10130), .Y(register__n1385) );
  HB1xp67_ASAP7_75t_R register___U4447 ( .A(register__n608), .Y(register__n12069) );
  HB1xp67_ASAP7_75t_R register___U4448 ( .A(register__n5045), .Y(register__n4576) );
  HB1xp67_ASAP7_75t_R register___U4449 ( .A(register__n5045), .Y(register__n4577) );
  HB1xp67_ASAP7_75t_R register___U4450 ( .A(register__n12585), .Y(register__n4426) );
  AO22x1_ASAP7_75t_R register___U4451 ( .A1(register__n9774), .A2(register__n387), .B1(register__n10275), .B2(register__net120912), .Y(register__n10691) );
  INVxp67_ASAP7_75t_R register___U4452 ( .A(register__n4521), .Y(register__n7038) );
  HB1xp67_ASAP7_75t_R register___U4453 ( .A(register__n4522), .Y(register__n4521) );
  HB1xp67_ASAP7_75t_R register___U4454 ( .A(register__n4919), .Y(register__n4918) );
  AND2x2_ASAP7_75t_R register___U4455 ( .A(register__n11601), .B(register__n11600), .Y(register__n1386) );
  NAND2xp33_ASAP7_75t_R register___U4456 ( .A(register__n1388), .B(register__n2117), .Y(register__n2308) );
  CKINVDCx20_ASAP7_75t_R register___U4457 ( .A(register__net94160), .Y(register__n1388) );
  INVxp67_ASAP7_75t_R register___U4458 ( .A(register__n3581), .Y(register__n5380) );
  NOR2xp67_ASAP7_75t_R register___U4459 ( .A(register__n1171), .B(register__n2695), .Y(register__n2697) );
  HB1xp67_ASAP7_75t_R register___U4460 ( .A(register__net105198), .Y(register__net64784) );
  INVx1_ASAP7_75t_R register___U4461 ( .A(register__n13260), .Y(register__n1389) );
  HB1xp67_ASAP7_75t_R register___U4462 ( .A(register__n12980), .Y(register__n5273) );
  NAND2xp33_ASAP7_75t_R register___U4463 ( .A(register__net90233), .B(register__n1867), .Y(register__n1390) );
  NAND2xp33_ASAP7_75t_R register___U4464 ( .A(register__net98195), .B(register__n1355), .Y(register__n1391) );
  NAND2xp33_ASAP7_75t_R register___U4465 ( .A(register__n1390), .B(register__n1391), .Y(register__n11088) );
  BUFx6f_ASAP7_75t_R register___U4466 ( .A(register__net109902), .Y(register__net90233) );
  HB1xp67_ASAP7_75t_R register___U4467 ( .A(register__net89017), .Y(register__net98195) );
  INVx6_ASAP7_75t_R register___U4468 ( .A(register__net64046), .Y(register__net64012) );
  INVxp33_ASAP7_75t_R register___U4469 ( .A(register__net64034), .Y(register__net64000) );
  INVx2_ASAP7_75t_R register___U4470 ( .A(register__n3159), .Y(register__n1544) );
  HB1xp67_ASAP7_75t_R register___U4471 ( .A(register__n5969), .Y(register__n5968) );
  INVx1_ASAP7_75t_R register___U4472 ( .A(register__n13246), .Y(register__n1392) );
  AOI22xp33_ASAP7_75t_R register___U4473 ( .A1(register__n12356), .A2(register__n11872), .B1(register__n1393), .B2(
        n1708), .Y(register__n13248) );
  INVx2_ASAP7_75t_R register___U4474 ( .A(register__n12356), .Y(register__n12338) );
  HB1xp67_ASAP7_75t_R register___U4475 ( .A(register__net64818), .Y(register__net64798) );
  INVxp67_ASAP7_75t_R register___U4476 ( .A(register__n11578), .Y(register__n4640) );
  AOI22xp33_ASAP7_75t_R register___U4477 ( .A1(register__n12133), .A2(register__n1112), .B1(register__n1394), .B2(register__n1701), .Y(register__n13252) );
  CKINVDCx20_ASAP7_75t_R register___U4478 ( .A(register__n10227), .Y(register__n1394) );
  INVxp67_ASAP7_75t_R register___U4479 ( .A(register__n4397), .Y(register__n7620) );
  AO22x2_ASAP7_75t_R register___U4480 ( .A1(register__net64056), .A2(register__n11731), .B1(register__n2708), .B2(register__n2021), .Y(register__n1395) );
  INVx1_ASAP7_75t_R register___U4481 ( .A(register__net64056), .Y(register__net63992) );
  CKINVDCx14_ASAP7_75t_R register___U4482 ( .A(register__n11731), .Y(register__n2021) );
  INVx1_ASAP7_75t_R register___U4483 ( .A(register__n13239), .Y(register__n1396) );
  INVxp67_ASAP7_75t_R register___U4484 ( .A(register__n6506), .Y(register__n8660) );
  HB1xp67_ASAP7_75t_R register___U4485 ( .A(register__n11069), .Y(register__n3498) );
  INVxp67_ASAP7_75t_R register___U4486 ( .A(register__net124480), .Y(register__net111717) );
  BUFx10_ASAP7_75t_R register___U4487 ( .A(register__net122410), .Y(register__net140639) );
  AND4x1_ASAP7_75t_R register___U4488 ( .A(register__n7072), .B(register__n5722), .C(register__n7071), .D(register__n3494), .Y(
        n10549) );
  HB1xp67_ASAP7_75t_R register___U4489 ( .A(register__n2872), .Y(register__n2871) );
  HB1xp67_ASAP7_75t_R register___U4490 ( .A(register__n11426), .Y(register__n2872) );
  AO22x1_ASAP7_75t_R register___U4491 ( .A1(register__n9270), .A2(register__C6422_net60408), .B1(register__n10193), 
        .B2(register__n838), .Y(register__n10790) );
  INVxp33_ASAP7_75t_R register___U4492 ( .A(register__n1951), .Y(register__n1813) );
  INVxp33_ASAP7_75t_R register___U4493 ( .A(register__n1813), .Y(register__n1814) );
  INVxp33_ASAP7_75t_R register___U4494 ( .A(register__n3711), .Y(register__n1817) );
  INVxp33_ASAP7_75t_R register___U4495 ( .A(register__n1817), .Y(register__n1818) );
  INVxp33_ASAP7_75t_R register___U4496 ( .A(register__n3709), .Y(register__n1821) );
  HB1xp67_ASAP7_75t_R register___U4497 ( .A(register__n11610), .Y(register__n4564) );
  INVxp67_ASAP7_75t_R register___U4498 ( .A(register__n4212), .Y(register__n7288) );
  HB1xp67_ASAP7_75t_R register___U4499 ( .A(register__n4213), .Y(register__n4212) );
  HB1xp67_ASAP7_75t_R register___U4500 ( .A(register__n12819), .Y(register__n3784) );
  INVxp67_ASAP7_75t_R register___U4501 ( .A(register__n13230), .Y(register__n4857) );
  HB1xp67_ASAP7_75t_R register___U4502 ( .A(register__n4398), .Y(register__n4397) );
  CKINVDCx20_ASAP7_75t_R register___U4503 ( .A(register__n9345), .Y(register__n1397) );
  INVx13_ASAP7_75t_R register___U4504 ( .A(register__n9327), .Y(register__n1399) );
  BUFx4f_ASAP7_75t_R register___U4505 ( .A(register__net64710), .Y(register__net64718) );
  INVx2_ASAP7_75t_R register___U4506 ( .A(register__net62858), .Y(register__net62826) );
  INVx1_ASAP7_75t_R register___U4507 ( .A(register__n12883), .Y(register__n1400) );
  HB1xp67_ASAP7_75t_R register___U4508 ( .A(register__n6507), .Y(register__n6506) );
  HB1xp67_ASAP7_75t_R register___U4509 ( .A(register__n3582), .Y(register__n3581) );
  INVxp67_ASAP7_75t_R register___U4510 ( .A(register__n12856), .Y(register__n8673) );
  INVxp67_ASAP7_75t_R register___U4511 ( .A(register__n3400), .Y(register__n5723) );
  HB1xp67_ASAP7_75t_R register___U4512 ( .A(register__n3401), .Y(register__n3400) );
  AO22x1_ASAP7_75t_R register___U4513 ( .A1(register__n9258), .A2(register__net122599), .B1(register__n9995), .B2(
        C6423_net68766), .Y(register__n11231) );
  BUFx2_ASAP7_75t_R register___U4514 ( .A(register__n2899), .Y(register__n2898) );
  INVxp67_ASAP7_75t_R register___U4515 ( .A(register__n13252), .Y(register__n7628) );
  BUFx3_ASAP7_75t_R register___U4516 ( .A(register__n3560), .Y(register__n11748) );
  HB1xp67_ASAP7_75t_R register___U4517 ( .A(register__n2886), .Y(register__n3436) );
  BUFx12f_ASAP7_75t_R register___U4518 ( .A(register__n11869), .Y(register__n2855) );
  HB1xp67_ASAP7_75t_R register___U4519 ( .A(register__n11748), .Y(register__n11749) );
  HB1xp67_ASAP7_75t_R register___U4520 ( .A(register__n11747), .Y(register__n3297) );
  BUFx12f_ASAP7_75t_R register___U4521 ( .A(register__n2855), .Y(register__n3561) );
  CKINVDCx10_ASAP7_75t_R register___U4522 ( .A(register__n3561), .Y(register__n2851) );
  INVx2_ASAP7_75t_R register___U4523 ( .A(register__n2835), .Y(register__n2834) );
  CKINVDCx20_ASAP7_75t_R register___U4524 ( .A(register__n7556), .Y(register__n1402) );
  AO22x1_ASAP7_75t_R register___U4525 ( .A1(register__n9895), .A2(register__net110414), .B1(register__n10153), .B2(
        net117889), .Y(register__n11674) );
  INVxp67_ASAP7_75t_R register___U4526 ( .A(register__n3962), .Y(register__n5906) );
  AO22x1_ASAP7_75t_R register___U4527 ( .A1(register__n9585), .A2(register__n1105), .B1(register__n10006), .B2(register__n285), 
        .Y(register__n11445) );
  INVxp67_ASAP7_75t_R register___U4528 ( .A(register__n6254), .Y(register__n6991) );
  BUFx6f_ASAP7_75t_R register___U4529 ( .A(register__n12504), .Y(register__n11913) );
  BUFx12f_ASAP7_75t_R register___U4530 ( .A(register__net145523), .Y(register__net145773) );
  HB1xp67_ASAP7_75t_R register___U4531 ( .A(register__n12855), .Y(register__n5007) );
  HB1xp67_ASAP7_75t_R register___U4532 ( .A(register__n11238), .Y(register__n2899) );
  BUFx6f_ASAP7_75t_R register___U4533 ( .A(register__n4818), .Y(register__n3603) );
  HB1xp67_ASAP7_75t_R register___U4534 ( .A(register__n12787), .Y(register__n4213) );
  HB1xp67_ASAP7_75t_R register___U4535 ( .A(register__n3963), .Y(register__n3962) );
  HB1xp67_ASAP7_75t_R register___U4536 ( .A(register__n4334), .Y(register__n4919) );
  INVx1_ASAP7_75t_R register___U4537 ( .A(register__n13321), .Y(register__n1404) );
  HB1xp67_ASAP7_75t_R register___U4538 ( .A(register__net124481), .Y(register__net124480) );
  INVx1_ASAP7_75t_R register___U4539 ( .A(register__n12573), .Y(register__n1405) );
  HB1xp67_ASAP7_75t_R register___U4540 ( .A(register__n549), .Y(register__n2828) );
  HB1xp67_ASAP7_75t_R register___U4541 ( .A(register__n13248), .Y(register__n4398) );
  HB1xp67_ASAP7_75t_R register___U4542 ( .A(register__n12816), .Y(register__n6507) );
  AO22x1_ASAP7_75t_R register___U4543 ( .A1(register__n9595), .A2(register__net93569), .B1(register__n10016), .B2(register__n284), 
        .Y(register__n11172) );
  INVxp33_ASAP7_75t_R register___U4544 ( .A(register__n7633), .Y(register__n1811) );
  HB1xp67_ASAP7_75t_R register___U4545 ( .A(register__n6255), .Y(register__n6254) );
  HB1xp67_ASAP7_75t_R register___U4546 ( .A(register__n13053), .Y(register__n5102) );
  AOI22x1_ASAP7_75t_R register___U4547 ( .A1(register__net63280), .A2(register__n904), .B1(register__n1756), .B2(register__n895), 
        .Y(register__n13044) );
  INVx1_ASAP7_75t_R register___U4548 ( .A(register__n12564), .Y(register__n1406) );
  INVxp33_ASAP7_75t_R register___U4549 ( .A(register__n3405), .Y(register__n6441) );
  INVxp67_ASAP7_75t_R register___U4550 ( .A(register__n3924), .Y(register__n5540) );
  HB1xp67_ASAP7_75t_R register___U4551 ( .A(register__n12925), .Y(register__n3963) );
  HB1xp67_ASAP7_75t_R register___U4552 ( .A(register__n13245), .Y(register__n6255) );
  INVxp67_ASAP7_75t_R register___U4553 ( .A(register__n13071), .Y(register__n8605) );
  INVx2_ASAP7_75t_R register___U4554 ( .A(register__n3120), .Y(register__n1545) );
  CKINVDCx20_ASAP7_75t_R register___U4555 ( .A(register__n9909), .Y(register__n1410) );
  INVx1_ASAP7_75t_R register___U4556 ( .A(register__n5721), .Y(register__n1414) );
  BUFx3_ASAP7_75t_R register___U4557 ( .A(register__n11834), .Y(register__n11832) );
  BUFx3_ASAP7_75t_R register___U4558 ( .A(register__n2984), .Y(register__n2961) );
  INVx6_ASAP7_75t_R register___U4559 ( .A(register__net64734), .Y(register__net144805) );
  BUFx12f_ASAP7_75t_R register___U4560 ( .A(register__net144805), .Y(register__net64732) );
  BUFx12f_ASAP7_75t_R register___U4561 ( .A(register__n11766), .Y(register__n1411) );
  HB1xp67_ASAP7_75t_R register___U4562 ( .A(register__n6441), .Y(register__n3404) );
  BUFx4f_ASAP7_75t_R register___U4563 ( .A(register__n5473), .Y(register__n5472) );
  HB1xp67_ASAP7_75t_R register___U4564 ( .A(register__n6782), .Y(register__n6781) );
  INVx1_ASAP7_75t_R register___U4565 ( .A(register__n11031), .Y(register__n1421) );
  BUFx6f_ASAP7_75t_R register___U4566 ( .A(register__n75), .Y(register__net108158) );
  BUFx6f_ASAP7_75t_R register___U4567 ( .A(register__net108158), .Y(register__C6422_net70602) );
  INVx1_ASAP7_75t_R register___U4568 ( .A(register__n13062), .Y(register__n1423) );
  AO22x1_ASAP7_75t_R register___U4569 ( .A1(register__n5443), .A2(register__n1417), .B1(register__n1759), .B2(register__n1415), 
        .Y(register__n1758) );
  INVx1_ASAP7_75t_R register___U4570 ( .A(register__n12716), .Y(register__n1424) );
  INVxp33_ASAP7_75t_R register___U4571 ( .A(register__n3071), .Y(register__n2139) );
  CKINVDCx20_ASAP7_75t_R register___U4572 ( .A(register__net90865), .Y(register__n1426) );
  AO22x1_ASAP7_75t_R register___U4573 ( .A1(register__n9290), .A2(register__n768), .B1(register__n9937), .B2(register__n75), .Y(
        n10630) );
  AO22x1_ASAP7_75t_R register___U4574 ( .A1(register__n9280), .A2(register__n768), .B1(register__n9933), .B2(register__n75), .Y(
        n10880) );
  AO22x1_ASAP7_75t_R register___U4575 ( .A1(register__net93853), .A2(register__C6422_net60408), .B1(register__net89793), 
        .B2(register__n835), .Y(register__n11001) );
  INVxp67_ASAP7_75t_R register___U4576 ( .A(register__n4013), .Y(register__n5948) );
  HB1xp67_ASAP7_75t_R register___U4577 ( .A(register__n4014), .Y(register__n4013) );
  AO22x1_ASAP7_75t_R register___U4578 ( .A1(register__n9836), .A2(register__net93569), .B1(register__n10253), .B2(
        C6423_net74857), .Y(register__n11598) );
  INVxp33_ASAP7_75t_R register___U4579 ( .A(register__n2970), .Y(register__n1595) );
  HB1xp67_ASAP7_75t_R register___U4580 ( .A(register__n3925), .Y(register__n3924) );
  AOI22xp33_ASAP7_75t_R register___U4581 ( .A1(register__n12099), .A2(register__n1695), .B1(register__n1427), .B2(register__n1710), .Y(register__n13255) );
  BUFx4f_ASAP7_75t_R register___U4582 ( .A(register__net64872), .Y(register__net64894) );
  INVx3_ASAP7_75t_R register___U4583 ( .A(register__net64894), .Y(register__net64858) );
  BUFx2_ASAP7_75t_R register___U4584 ( .A(register__n11366), .Y(register__n5916) );
  INVxp33_ASAP7_75t_R register___U4585 ( .A(register__n4851), .Y(register__n1848) );
  INVxp33_ASAP7_75t_R register___U4586 ( .A(register__n4851), .Y(register__n1849) );
  AOI22xp33_ASAP7_75t_R register___U4587 ( .A1(register__n9296), .A2(register__n77), .B1(register__n10446), .B2(register__n75), 
        .Y(register__n1429) );
  BUFx12f_ASAP7_75t_R register___U4588 ( .A(register__net62680), .Y(register__net144425) );
  CKINVDCx20_ASAP7_75t_R register___U4589 ( .A(register__n9413), .Y(register__n1430) );
  CKINVDCx5p33_ASAP7_75t_R register___U4590 ( .A(register__net141489), .Y(register__net64676) );
  BUFx6f_ASAP7_75t_R register___U4591 ( .A(register__net66306), .Y(register__net66308) );
  HB1xp67_ASAP7_75t_R register___U4592 ( .A(register__n10622), .Y(register__n4334) );
  AO22x1_ASAP7_75t_R register___U4593 ( .A1(register__n6670), .A2(register__n768), .B1(register__n10315), .B2(
        C6422_net60437), .Y(register__n10856) );
  HB1xp67_ASAP7_75t_R register___U4594 ( .A(register__n13094), .Y(register__n3925) );
  AO22x1_ASAP7_75t_R register___U4595 ( .A1(register__net93639), .A2(register__net117657), .B1(register__net96819), 
        .B2(register__n838), .Y(register__n10806) );
  INVxp67_ASAP7_75t_R register___U4596 ( .A(register__n2971), .Y(register__n3663) );
  BUFx3_ASAP7_75t_R register___U4597 ( .A(register__n11912), .Y(register__n7973) );
  HB1xp67_ASAP7_75t_R register___U4598 ( .A(register__n6253), .Y(register__n6252) );
  AO22x1_ASAP7_75t_R register___U4599 ( .A1(register__n9712), .A2(register__net131160), .B1(register__n10042), .B2(
        net120912), .Y(register__n10672) );
  NOR4xp75_ASAP7_75t_R register___U4600 ( .A(register__n11285), .B(register__n4101), .C(register__n11287), .D(register__n1433), 
        .Y(register__n11280) );
  HB1xp67_ASAP7_75t_R register___U4601 ( .A(register__n12691), .Y(register__n6253) );
  AOI22xp33_ASAP7_75t_R register___U4602 ( .A1(register__n6097), .A2(register__net106379), .B1(register__n10124), .B2(
        n2000), .Y(register__n1434) );
  INVx1_ASAP7_75t_R register___U4603 ( .A(register__n11615), .Y(register__n3591) );
  HB1xp67_ASAP7_75t_R register___U4604 ( .A(register__n2972), .Y(register__n2971) );
  INVx2_ASAP7_75t_R register___U4605 ( .A(register__n12264), .Y(register__n12252) );
  OAI22xp5_ASAP7_75t_R register___U4606 ( .A1(register__net66304), .A2(register__n7613), .B1(register__net64696), .B2(
        n1687), .Y(read_reg_data_2[7]) );
  INVxp67_ASAP7_75t_R register___U4607 ( .A(register__n13255), .Y(register__n7626) );
  INVx1_ASAP7_75t_R register___U4608 ( .A(register__n13259), .Y(register__n1436) );
  INVx2_ASAP7_75t_R register___U4609 ( .A(register__n2765), .Y(register__n1458) );
  HB1xp67_ASAP7_75t_R register___U4610 ( .A(register__n12991), .Y(register__n4149) );
  AOI22xp33_ASAP7_75t_R register___U4611 ( .A1(register__n9736), .A2(register__C6423_net61326), .B1(register__n9319), 
        .B2(register__n2001), .Y(register__n1437) );
  OA22x2_ASAP7_75t_R register___U4612 ( .A1(register__n1438), .A2(register__n2419), .B1(register__n1751), .B2(register__n277), 
        .Y(register__n1482) );
  CKINVDCx20_ASAP7_75t_R register___U4613 ( .A(register__n9573), .Y(register__n1438) );
  INVx13_ASAP7_75t_R register___U4614 ( .A(register__n9429), .Y(register__n1751) );
  HB1xp67_ASAP7_75t_R register___U4615 ( .A(register__n11002), .Y(register__n2839) );
  AO22x1_ASAP7_75t_R register___U4616 ( .A1(register__net96903), .A2(register__n375), .B1(register__net90093), .B2(
        C6422_net60401), .Y(register__n11002) );
  HB1xp67_ASAP7_75t_R register___U4617 ( .A(register__n12947), .Y(register__n4778) );
  HB1xp67_ASAP7_75t_R register___U4618 ( .A(register__n12364), .Y(register__n5348) );
  INVxp33_ASAP7_75t_R register___U4619 ( .A(register__n1441), .Y(register__n1453) );
  INVxp33_ASAP7_75t_R register___U4620 ( .A(register__n1441), .Y(register__n1454) );
  BUFx12f_ASAP7_75t_R register___U4621 ( .A(register__n12008), .Y(register__n12005) );
  AO22x1_ASAP7_75t_R register___U4622 ( .A1(register__n8343), .A2(register__C6423_net61318), .B1(register__n10020), 
        .B2(register__n1445), .Y(register__n11530) );
  HB1xp67_ASAP7_75t_R register___U4623 ( .A(register__net36421), .Y(register__net124481) );
  INVxp67_ASAP7_75t_R register___U4624 ( .A(register__n11666), .Y(register__n7271) );
  HB1xp67_ASAP7_75t_R register___U4625 ( .A(register__n4849), .Y(register__n4265) );
  INVx2_ASAP7_75t_R register___U4626 ( .A(register__n4265), .Y(register__n12153) );
  AO22x1_ASAP7_75t_R register___U4627 ( .A1(register__n9889), .A2(register__n413), .B1(register__n10313), .B2(register__net126601), .Y(register__n10849) );
  HB1xp67_ASAP7_75t_R register___U4628 ( .A(register__n4145), .Y(register__n4144) );
  AO22x1_ASAP7_75t_R register___U4629 ( .A1(register__n9292), .A2(register__net122579), .B1(register__n9939), .B2(
        net150888), .Y(register__n11216) );
  INVxp67_ASAP7_75t_R register___U4630 ( .A(register__n13058), .Y(register__n9183) );
  HB1xp67_ASAP7_75t_R register___U4631 ( .A(register__n13278), .Y(register__n2972) );
  HB1xp67_ASAP7_75t_R register___U4632 ( .A(register__n12796), .Y(register__n6782) );
  BUFx12_ASAP7_75t_R register___U4633 ( .A(register__net140298), .Y(register__net139861) );
  INVx1_ASAP7_75t_R register___U4634 ( .A(register__n12685), .Y(register__n1456) );
  INVx1_ASAP7_75t_R register___U4635 ( .A(register__n11483), .Y(register__n1457) );
  AO22x1_ASAP7_75t_R register___U4636 ( .A1(register__n8805), .A2(register__net124706), .B1(register__n7337), .B2(register__n2000), .Y(register__n11483) );
  AO22x1_ASAP7_75t_R register___U4637 ( .A1(register__n9587), .A2(register__net93569), .B1(register__n10008), .B2(
        C6423_net74857), .Y(register__n11339) );
  INVx1_ASAP7_75t_R register___U4638 ( .A(register__n10853), .Y(register__n1460) );
  AND2x2_ASAP7_75t_R register___U4639 ( .A(register__n10547), .B(register__n7670), .Y(register__n1461) );
  AO22x1_ASAP7_75t_R register___U4640 ( .A1(register__net93741), .A2(register__net122579), .B1(register__net90113), 
        .B2(register__net150884), .Y(register__n11294) );
  AO22x1_ASAP7_75t_R register___U4641 ( .A1(register__net93737), .A2(register__n931), .B1(register__net90109), .B2(
        net150889), .Y(register__n11275) );
  BUFx2_ASAP7_75t_R register___U4642 ( .A(register__n4248), .Y(register__n4247) );
  HB1xp67_ASAP7_75t_R register___U4643 ( .A(register__n12769), .Y(register__n4145) );
  AO22x1_ASAP7_75t_R register___U4644 ( .A1(register__net90761), .A2(register__net131160), .B1(register__net89845), 
        .B2(register__net120912), .Y(register__n11007) );
  AO22x1_ASAP7_75t_R register___U4645 ( .A1(register__n9832), .A2(register__net131160), .B1(register__n10128), .B2(
        net120912), .Y(register__n10988) );
  HB1xp67_ASAP7_75t_R register___U4646 ( .A(register__n12017), .Y(register__n12003) );
  HB1xp67_ASAP7_75t_R register___U4647 ( .A(register__n12017), .Y(register__n12002) );
  HB1xp67_ASAP7_75t_R register___U4648 ( .A(register__n12017), .Y(register__n12001) );
  HB1xp67_ASAP7_75t_R register___U4649 ( .A(register__n12017), .Y(register__n12006) );
  AOI21xp33_ASAP7_75t_R register___U4650 ( .A1(register__net93569), .A2(register__net90453), .B(register__n2494), .Y(
        n2514) );
  AO22x1_ASAP7_75t_R register___U4651 ( .A1(register__n9094), .A2(register__n38), .B1(register__n10165), .B2(
        C6422_net60443), .Y(register__n11030) );
  HB1xp67_ASAP7_75t_R register___U4652 ( .A(register__n3605), .Y(register__n1462) );
  HB1xp67_ASAP7_75t_R register___U4653 ( .A(register__n3605), .Y(register__n1463) );
  BUFx12f_ASAP7_75t_R register___U4654 ( .A(register__n12500), .Y(register__n3217) );
  BUFx6f_ASAP7_75t_R register___U4655 ( .A(register__n4177), .Y(register__n4632) );
  BUFx3_ASAP7_75t_R register___U4656 ( .A(register__n3261), .Y(register__n11807) );
  BUFx6f_ASAP7_75t_R register___U4657 ( .A(register__n4632), .Y(register__n5685) );
  HB1xp67_ASAP7_75t_R register___U4658 ( .A(register__n11807), .Y(register__n5356) );
  HB1xp67_ASAP7_75t_R register___U4659 ( .A(register__n3508), .Y(register__n3477) );
  HB1xp67_ASAP7_75t_R register___U4660 ( .A(register__n5685), .Y(register__n3413) );
  HB1xp67_ASAP7_75t_R register___U4661 ( .A(register__n5685), .Y(register__n3414) );
  HB1xp67_ASAP7_75t_R register___U4662 ( .A(register__n11891), .Y(register__n11805) );
  INVxp67_ASAP7_75t_R register___U4663 ( .A(register__n4907), .Y(register__n8263) );
  INVxp67_ASAP7_75t_R register___U4664 ( .A(register__n3055), .Y(register__n1464) );
  BUFx3_ASAP7_75t_R register___U4665 ( .A(register__n11912), .Y(register__n3472) );
  HB1xp67_ASAP7_75t_R register___U4666 ( .A(register__n5742), .Y(register__n9169) );
  HB1xp67_ASAP7_75t_R register___U4667 ( .A(register__n5743), .Y(register__n5742) );
  HB1xp67_ASAP7_75t_R register___U4668 ( .A(register__n12794), .Y(register__n4502) );
  HB1xp67_ASAP7_75t_R register___U4669 ( .A(register__n12793), .Y(register__n6249) );
  INVxp67_ASAP7_75t_R register___U4670 ( .A(register__n13136), .Y(register__n3562) );
  INVxp67_ASAP7_75t_R register___U4671 ( .A(register__n3367), .Y(register__n4647) );
  HB1xp67_ASAP7_75t_R register___U4672 ( .A(register__n3368), .Y(register__n3367) );
  INVx6_ASAP7_75t_R register___U4673 ( .A(register__net64374), .Y(register__net64342) );
  HB1xp67_ASAP7_75t_R register___U4674 ( .A(register__n10901), .Y(register__n4248) );
  AO22x1_ASAP7_75t_R register___U4675 ( .A1(register__n9054), .A2(register__n387), .B1(register__n8376), .B2(register__n326), .Y(
        n11115) );
  INVx1_ASAP7_75t_R register___U4676 ( .A(register__n11460), .Y(register__n1465) );
  BUFx6f_ASAP7_75t_R register___U4677 ( .A(register__n11767), .Y(register__n11766) );
  INVxp67_ASAP7_75t_R register___U4678 ( .A(register__n1758), .Y(register__n12994) );
  INVxp67_ASAP7_75t_R register___U4679 ( .A(register__n3771), .Y(register__n5901) );
  AO22x1_ASAP7_75t_R register___U4680 ( .A1(register__n1467), .A2(register__n1470), .B1(register__n1468), .B2(register__n1469), 
        .Y(read_reg_data_2[3]) );
  CKINVDCx20_ASAP7_75t_R register___U4681 ( .A(register__n12033), .Y(register__n1468) );
  CKINVDCx20_ASAP7_75t_R register___U4682 ( .A(register__n1687), .Y(register__n1469) );
  OAI22xp5_ASAP7_75t_R register___U4683 ( .A1(register__n1471), .A2(register__n11889), .B1(register__n10446), .B2(register__n7656), .Y(register__n2219) );
  BUFx2_ASAP7_75t_R register___U4684 ( .A(register__n4448), .Y(register__n4447) );
  INVx1_ASAP7_75t_R register___U4685 ( .A(register__n12478), .Y(register__n12462) );
  INVx1_ASAP7_75t_R register___U4686 ( .A(register__n11626), .Y(register__n1472) );
  HB1xp67_ASAP7_75t_R register___U4687 ( .A(register__n13386), .Y(register__n4014) );
  HB1xp67_ASAP7_75t_R register___U4688 ( .A(register__n3021), .Y(register__n1474) );
  OAI22xp33_ASAP7_75t_R register___U4689 ( .A1(register__n3644), .A2(register__n109), .B1(register__n9965), .B2(register__n5504), 
        .Y(register__n1475) );
  AND2x2_ASAP7_75t_R register___U4690 ( .A(register__n12495), .B(register__n12485), .Y(register__n12499) );
  BUFx6f_ASAP7_75t_R register___U4691 ( .A(register__n12499), .Y(register__n1774) );
  HB1xp67_ASAP7_75t_R register___U4692 ( .A(register__n5838), .Y(register__n3307) );
  BUFx6f_ASAP7_75t_R register___U4693 ( .A(register__n5660), .Y(register__n11886) );
  NOR2xp67_ASAP7_75t_R register___U4694 ( .A(register__n2307), .B(register__n1889), .Y(register__net36421) );
  INVx1_ASAP7_75t_R register___U4695 ( .A(register__n2308), .Y(register__n1889) );
  HB1xp67_ASAP7_75t_R register___U4696 ( .A(register__n4908), .Y(register__n4907) );
  BUFx12f_ASAP7_75t_R register___U4697 ( .A(register__net141466), .Y(register__net142763) );
  HB1xp67_ASAP7_75t_R register___U4698 ( .A(register__n12837), .Y(register__n4664) );
  INVxp67_ASAP7_75t_R register___U4699 ( .A(register__n13116), .Y(register__n8556) );
  AND2x2_ASAP7_75t_R register___U4700 ( .A(register__n566), .B(register__n8251), .Y(register__n1477) );
  AND4x1_ASAP7_75t_R register___U4701 ( .A(register__n11473), .B(register__n8284), .C(register__n11474), .D(register__n11472), 
        .Y(register__n8584) );
  AO22x1_ASAP7_75t_R register___U4702 ( .A1(register__n6916), .A2(register__n768), .B1(register__n9382), .B2(register__n75), .Y(
        n10947) );
  NOR4xp75_ASAP7_75t_R register___U4703 ( .A(register__n5621), .B(register__n1478), .C(register__n1479), .D(register__n4910), .Y(
        n11408) );
  BUFx6f_ASAP7_75t_R register___U4704 ( .A(register__net140270), .Y(register__net64380) );
  AO22x1_ASAP7_75t_R register___U4705 ( .A1(register__n9724), .A2(register__n387), .B1(register__n10175), .B2(register__net120912), .Y(register__n10853) );
  AO22x1_ASAP7_75t_R register___U4706 ( .A1(register__net93717), .A2(register__n925), .B1(register__net89041), .B2(
        net150882), .Y(register__n11614) );
  AO22x1_ASAP7_75t_R register___U4707 ( .A1(register__n6656), .A2(register__net122579), .B1(register__n10261), .B2(
        net121558), .Y(register__n11597) );
  AO22x1_ASAP7_75t_R register___U4708 ( .A1(register__n5175), .A2(register__n1106), .B1(register__n6050), .B2(register__n285), 
        .Y(register__n11238) );
  HB1xp67_ASAP7_75t_R register___U4709 ( .A(register__n4650), .Y(register__n12210) );
  HB1xp67_ASAP7_75t_R register___U4710 ( .A(register__n11117), .Y(register__n4908) );
  HB1xp67_ASAP7_75t_R register___U4711 ( .A(register__n6404), .Y(register__n4649) );
  HB1xp67_ASAP7_75t_R register___U4712 ( .A(register__n3772), .Y(register__n3771) );
  BUFx2_ASAP7_75t_R register___U4713 ( .A(register__n4623), .Y(register__n8257) );
  AND3x2_ASAP7_75t_R register___U4714 ( .A(register__n11721), .B(register__n731), .C(register__n5441), .Y(register__n11720) );
  HB1xp67_ASAP7_75t_R register___U4715 ( .A(register__n4624), .Y(register__n4623) );
  OAI22xp5_ASAP7_75t_R register___U4716 ( .A1(register__net66312), .A2(register__n8584), .B1(register__n12266), .B2(
        n1687), .Y(read_reg_data_2[18]) );
  INVx1_ASAP7_75t_R register___U4717 ( .A(register__n12550), .Y(register__n1485) );
  BUFx6f_ASAP7_75t_R register___U4718 ( .A(register__n4604), .Y(register__n4603) );
  HB1xp67_ASAP7_75t_R register___U4719 ( .A(register__n12541), .Y(register__n4299) );
  BUFx6f_ASAP7_75t_R register___U4720 ( .A(register__n11839), .Y(register__n11841) );
  BUFx2_ASAP7_75t_R register___U4721 ( .A(register__n3361), .Y(register__n5050) );
  CKINVDCx10_ASAP7_75t_R register___U4722 ( .A(register__net142571), .Y(register__net117320) );
  HB1xp67_ASAP7_75t_R register___U4723 ( .A(register__net63390), .Y(register__net63362) );
  HB1xp67_ASAP7_75t_R register___U4724 ( .A(register__net63390), .Y(register__net63366) );
  HB1xp67_ASAP7_75t_R register___U4725 ( .A(register__n11688), .Y(register__n4624) );
  INVx6_ASAP7_75t_R register___U4726 ( .A(register__net62856), .Y(register__net62824) );
  BUFx12f_ASAP7_75t_R register___U4727 ( .A(register__net121482), .Y(register__net62856) );
  INVx2_ASAP7_75t_R register___U4728 ( .A(register__n4716), .Y(register__n6711) );
  HB1xp67_ASAP7_75t_R register___U4729 ( .A(register__n12904), .Y(register__n3165) );
  INVx1_ASAP7_75t_R register___U4730 ( .A(register__n13054), .Y(register__n1486) );
  AO22x1_ASAP7_75t_R register___U4731 ( .A1(register__n6910), .A2(register__n923), .B1(register__n9941), .B2(register__n1898), 
        .Y(register__n11171) );
  CKINVDCx20_ASAP7_75t_R register___U4732 ( .A(register__n10018), .Y(register__n1488) );
  HB1xp67_ASAP7_75t_R register___U4733 ( .A(register__n13272), .Y(register__n3405) );
  INVxp67_ASAP7_75t_R register___U4734 ( .A(register__n5775), .Y(register__n7625) );
  AO22x1_ASAP7_75t_R register___U4735 ( .A1(register__n9347), .A2(register__net128121), .B1(register__n9365), .B2(register__n2000), .Y(register__n11626) );
  HB1xp67_ASAP7_75t_R register___U4736 ( .A(register__n12998), .Y(register__n3368) );
  CKINVDCx10_ASAP7_75t_R register___U4737 ( .A(register__net144944), .Y(register__net142571) );
  CKINVDCx20_ASAP7_75t_R register___U4738 ( .A(register__n6610), .Y(register__n1491) );
  NAND2xp33_ASAP7_75t_R register___U4739 ( .A(register__n9623), .B(register__net110414), .Y(register__n1492) );
  NAND2xp33_ASAP7_75t_R register___U4740 ( .A(register__n1492), .B(register__n1493), .Y(register__n11536) );
  AND2x2_ASAP7_75t_R register___U4741 ( .A(register__n11519), .B(register__n376), .Y(register__n1494) );
  AND3x1_ASAP7_75t_R register___U4742 ( .A(register__n1494), .B(register__n11517), .C(register__n11518), .Y(register__n6162) );
  HB1xp67_ASAP7_75t_R register___U4743 ( .A(register__n10086), .Y(register__n7486) );
  INVxp67_ASAP7_75t_R register___U4744 ( .A(register__n10544), .Y(register__n7878) );
  HB1xp67_ASAP7_75t_R register___U4745 ( .A(register__n11533), .Y(register__n4311) );
  OAI22xp5_ASAP7_75t_R register___U4746 ( .A1(register__net66312), .A2(register__n4178), .B1(register__n12294), .B2(
        n1687), .Y(read_reg_data_2[19]) );
  AOI21xp33_ASAP7_75t_R register___U4747 ( .A1(register__C6423_net68764), .A2(register__net89969), .B(register__n2415), 
        .Y(register__n2438) );
  AO22x1_ASAP7_75t_R register___U4748 ( .A1(register__n9415), .A2(register__net138603), .B1(register__n7215), .B2(
        net125803), .Y(register__n11591) );
  INVxp67_ASAP7_75t_R register___U4749 ( .A(register__n12838), .Y(register__n8676) );
  INVx4_ASAP7_75t_R register___U4750 ( .A(register__net64698), .Y(register__net64664) );
  INVx1_ASAP7_75t_R register___U4751 ( .A(register__n13264), .Y(register__n1497) );
  OAI22xp33_ASAP7_75t_R register___U4752 ( .A1(register__n12402), .A2(register__n109), .B1(register__n10114), .B2(
        n11887), .Y(register__n1498) );
  INVx1_ASAP7_75t_R register___U4753 ( .A(register__n12863), .Y(register__n1499) );
  AO22x1_ASAP7_75t_R register___U4754 ( .A1(register__n9621), .A2(register__net110414), .B1(register__n10076), .B2(
        net125797), .Y(register__n11576) );
  HB1xp67_ASAP7_75t_R register___U4755 ( .A(register__n12824), .Y(register__n3521) );
  HB1xp67_ASAP7_75t_R register___U4756 ( .A(register__n12807), .Y(register__n5406) );
  HB1xp67_ASAP7_75t_R register___U4757 ( .A(register__n3612), .Y(register__n3611) );
  HB1xp67_ASAP7_75t_R register___U4758 ( .A(register__n12815), .Y(register__n3612) );
  INVxp67_ASAP7_75t_R register___U4759 ( .A(register__n4082), .Y(register__n4183) );
  HB1xp67_ASAP7_75t_R register___U4760 ( .A(register__n12935), .Y(register__n4782) );
  BUFx6f_ASAP7_75t_R register___U4761 ( .A(register__n3374), .Y(register__n4727) );
  BUFx12f_ASAP7_75t_R register___U4762 ( .A(register__net117320), .Y(register__net64374) );
  AO22x1_ASAP7_75t_R register___U4763 ( .A1(register__n6911), .A2(register__n77), .B1(register__n9941), .B2(register__n75), .Y(
        n10544) );
  INVxp67_ASAP7_75t_R register___U4764 ( .A(register__n2948), .Y(register__n3592) );
  AO22x1_ASAP7_75t_R register___U4765 ( .A1(register__net96843), .A2(register__net126316), .B1(register__net91583), 
        .B2(register__net123880), .Y(register__n11089) );
  INVx2_ASAP7_75t_R register___U4766 ( .A(register__n11693), .Y(register__n6709) );
  HB1xp67_ASAP7_75t_R register___U4767 ( .A(register__n5776), .Y(register__n5775) );
  INVx1_ASAP7_75t_R register___U4768 ( .A(register__n11266), .Y(register__n1502) );
  INVxp67_ASAP7_75t_R register___U4769 ( .A(register__n7352), .Y(register__n8681) );
  INVxp67_ASAP7_75t_R register___U4770 ( .A(register__n3857), .Y(register__n5370) );
  AO22x1_ASAP7_75t_R register___U4771 ( .A1(register__n9796), .A2(register__net126316), .B1(register__n10116), .B2(
        net123880), .Y(register__n11113) );
  BUFx3_ASAP7_75t_R register___U4772 ( .A(register__n11047), .Y(register__n7305) );
  INVxp67_ASAP7_75t_R register___U4773 ( .A(register__n4413), .Y(register__n8683) );
  HB1xp67_ASAP7_75t_R register___U4774 ( .A(register__n12828), .Y(register__n3656) );
  HB1xp67_ASAP7_75t_R register___U4775 ( .A(register__n6266), .Y(register__n6059) );
  INVx6_ASAP7_75t_R register___U4776 ( .A(register__net64062), .Y(register__net120674) );
  HB1xp67_ASAP7_75t_R register___U4777 ( .A(register__net120674), .Y(register__net129902) );
  BUFx12f_ASAP7_75t_R register___U4778 ( .A(register__net142960), .Y(register__net144944) );
  INVxp67_ASAP7_75t_R register___U4779 ( .A(register__n4417), .Y(register__n9164) );
  HB1xp67_ASAP7_75t_R register___U4780 ( .A(register__n4418), .Y(register__n4417) );
  INVxp67_ASAP7_75t_R register___U4781 ( .A(register__n4541), .Y(register__n8624) );
  HB1xp67_ASAP7_75t_R register___U4782 ( .A(register__n4542), .Y(register__n4541) );
  INVx1_ASAP7_75t_R register___U4783 ( .A(register__n11538), .Y(register__n1504) );
  HB1xp67_ASAP7_75t_R register___U4784 ( .A(register__n4083), .Y(register__n4082) );
  INVxp67_ASAP7_75t_R register___U4785 ( .A(register__n4477), .Y(register__n7921) );
  AO22x1_ASAP7_75t_R register___U4786 ( .A1(register__net114452), .A2(register__net113802), .B1(register__net91563), 
        .B2(register__C6423_net68766), .Y(register__n11288) );
  INVxp67_ASAP7_75t_R register___U4787 ( .A(register__n5312), .Y(register__n5912) );
  HB1xp67_ASAP7_75t_R register___U4788 ( .A(register__n5313), .Y(register__n5312) );
  BUFx6f_ASAP7_75t_R register___U4789 ( .A(register__n7258), .Y(register__n12447) );
  INVx1_ASAP7_75t_R register___U4790 ( .A(register__n11167), .Y(register__n1505) );
  HB1xp67_ASAP7_75t_R register___U4791 ( .A(register__n3551), .Y(register__n3550) );
  INVx1_ASAP7_75t_R register___U4792 ( .A(register__n11290), .Y(register__n1506) );
  HB1xp67_ASAP7_75t_R register___U4793 ( .A(register__n2949), .Y(register__n2948) );
  HB1xp67_ASAP7_75t_R register___U4794 ( .A(register__n3858), .Y(register__n3857) );
  NAND3xp33_ASAP7_75t_R register___U4795 ( .A(register__n12507), .B(register__n7679), .C(register__n7678), .Y(register__n1507) );
  CKINVDCx10_ASAP7_75t_R register___U4796 ( .A(register__net63198), .Y(register__net63166) );
  AO22x1_ASAP7_75t_R register___U4797 ( .A1(register__net91105), .A2(register__net106379), .B1(register__net89777), 
        .B2(register__n2000), .Y(register__n11285) );
  HB1xp67_ASAP7_75t_R register___U4798 ( .A(register__n11648), .Y(register__n5313) );
  AO22x1_ASAP7_75t_R register___U4799 ( .A1(register__n8809), .A2(register__net126316), .B1(register__n8353), .B2(
        net123880), .Y(register__n11047) );
  INVx1_ASAP7_75t_R register___U4800 ( .A(register__n11313), .Y(register__n1508) );
  HB1xp67_ASAP7_75t_R register___U4801 ( .A(register__n11311), .Y(register__n4336) );
  AO22x1_ASAP7_75t_R register___U4802 ( .A1(register__n9413), .A2(register__net125426), .B1(register__n10181), .B2(register__n162), .Y(register__n11311) );
  AO22x1_ASAP7_75t_R register___U4803 ( .A1(register__net93837), .A2(register__net124706), .B1(register__net89773), 
        .B2(register__n2001), .Y(register__n11266) );
  HB1xp67_ASAP7_75t_R register___U4804 ( .A(register__n2929), .Y(register__n4974) );
  HB1xp67_ASAP7_75t_R register___U4805 ( .A(register__n4478), .Y(register__n4477) );
  HB1xp67_ASAP7_75t_R register___U4806 ( .A(register__n7322), .Y(register__n4337) );
  AO22x1_ASAP7_75t_R register___U4807 ( .A1(register__n7515), .A2(register__C6423_net61318), .B1(register__n6629), .B2(
        n1447), .Y(register__n11310) );
  INVxp67_ASAP7_75t_R register___U4808 ( .A(register__n4172), .Y(register__n7058) );
  INVxp67_ASAP7_75t_R register___U4809 ( .A(register__n12693), .Y(register__n6683) );
  AND2x2_ASAP7_75t_R register___U4810 ( .A(register__n12485), .B(register__n12503), .Y(register__n6139) );
  BUFx4f_ASAP7_75t_R register___U4811 ( .A(register__n11903), .Y(register__n3756) );
  CKINVDCx6p67_ASAP7_75t_R register___U4812 ( .A(register__n4267), .Y(register__n4268) );
  BUFx6f_ASAP7_75t_R register___U4813 ( .A(register__n3756), .Y(register__n3547) );
  INVx1_ASAP7_75t_R register___U4814 ( .A(register__n11900), .Y(register__n5047) );
  BUFx6f_ASAP7_75t_R register___U4815 ( .A(register__n3547), .Y(register__n3327) );
  BUFx3_ASAP7_75t_R register___U4816 ( .A(register__n3547), .Y(register__n3328) );
  BUFx6f_ASAP7_75t_R register___U4817 ( .A(register__n3327), .Y(register__n11901) );
  BUFx6f_ASAP7_75t_R register___U4818 ( .A(register__n11824), .Y(register__n3152) );
  BUFx6f_ASAP7_75t_R register___U4819 ( .A(register__n11824), .Y(register__n3153) );
  BUFx3_ASAP7_75t_R register___U4820 ( .A(register__n11901), .Y(register__n5184) );
  BUFx3_ASAP7_75t_R register___U4821 ( .A(register__n11901), .Y(register__n11821) );
  BUFx3_ASAP7_75t_R register___U4822 ( .A(register__n3480), .Y(register__n3385) );
  BUFx3_ASAP7_75t_R register___U4823 ( .A(register__n3480), .Y(register__n3479) );
  HB1xp67_ASAP7_75t_R register___U4824 ( .A(register__n3153), .Y(register__n11823) );
  CKINVDCx20_ASAP7_75t_R register___U4825 ( .A(register__n11820), .Y(register__n4267) );
  CKINVDCx8_ASAP7_75t_R register___U4826 ( .A(register__n4268), .Y(register__n11900) );
  BUFx12f_ASAP7_75t_R register___U4827 ( .A(register__net140686), .Y(register__net63198) );
  INVxp67_ASAP7_75t_R register___U4828 ( .A(register__C6423_net68930), .Y(register__n_cell_125217_net175396)
         );
  HB1xp67_ASAP7_75t_R register___U4829 ( .A(register__n11570), .Y(register__n4478) );
  BUFx6f_ASAP7_75t_R register___U4830 ( .A(register__n1861), .Y(register__n11764) );
  INVxp67_ASAP7_75t_R register___U4831 ( .A(register__n3125), .Y(register__n5382) );
  HB1xp67_ASAP7_75t_R register___U4832 ( .A(register__n3126), .Y(register__n3125) );
  AO22x1_ASAP7_75t_R register___U4833 ( .A1(register__n9840), .A2(register__n128), .B1(register__n8170), .B2(register__n1445), 
        .Y(register__n11648) );
  HB1xp67_ASAP7_75t_R register___U4834 ( .A(register__n2930), .Y(register__n2929) );
  INVxp67_ASAP7_75t_R register___U4835 ( .A(register__n10816), .Y(register__n7915) );
  HB1xp67_ASAP7_75t_R register___U4836 ( .A(register__n11716), .Y(register__n4172) );
  AOI21xp33_ASAP7_75t_R register___U4837 ( .A1(register__net94399), .A2(register__net90093), .B(register__n2417), .Y(
        n2441) );
  AO22x1_ASAP7_75t_R register___U4838 ( .A1(register__n8763), .A2(register__net125170), .B1(register__n9359), .B2(register__n515), 
        .Y(register__n11185) );
  AO22x1_ASAP7_75t_R register___U4839 ( .A1(register__n9845), .A2(register__net125170), .B1(register__n6649), .B2(register__n515), 
        .Y(register__n11589) );
  AO22x1_ASAP7_75t_R register___U4840 ( .A1(register__net90537), .A2(register__net125170), .B1(register__net89045), 
        .B2(register__n235), .Y(register__n11607) );
  HB1xp67_ASAP7_75t_R register___U4841 ( .A(register__n4608), .Y(register__n4607) );
  HB1xp67_ASAP7_75t_R register___U4842 ( .A(register__n11251), .Y(register__n4608) );
  AO22x1_ASAP7_75t_R register___U4843 ( .A1(register__n9329), .A2(register__n1035), .B1(register__n7467), .B2(register__n2000), 
        .Y(register__n11184) );
  AO22x1_ASAP7_75t_R register___U4844 ( .A1(register__n9577), .A2(register__C6423_net61326), .B1(register__n10062), 
        .B2(register__n2001), .Y(register__n11162) );
  AO22x1_ASAP7_75t_R register___U4845 ( .A1(register__n9810), .A2(register__net125170), .B1(register__n10335), .B2(register__n235), .Y(register__n11667) );
  AND4x2_ASAP7_75t_R register___U4846 ( .A(register__n4740), .B(register__n7073), .C(register__n5912), .D(register__n2252), .Y(
        n11640) );
  AO22x1_ASAP7_75t_R register___U4847 ( .A1(register__n9587), .A2(register__n1771), .B1(register__n10008), .B2(
        net126625), .Y(register__n10676) );
  HB1xp67_ASAP7_75t_R register___U4848 ( .A(register__n11310), .Y(register__n5743) );
  INVxp67_ASAP7_75t_R register___U4849 ( .A(register__n5276), .Y(register__n6999) );
  INVx1_ASAP7_75t_R register___U4850 ( .A(register__n4911), .Y(register__n7272) );
  INVx1_ASAP7_75t_R register___U4851 ( .A(register__n11700), .Y(register__n2275) );
  AO22x1_ASAP7_75t_R register___U4852 ( .A1(register__n9640), .A2(register__net125170), .B1(register__n9951), .B2(register__n515), 
        .Y(register__n11163) );
  AO22x1_ASAP7_75t_R register___U4853 ( .A1(register__n9873), .A2(register__net125170), .B1(register__n10287), .B2(register__n515), .Y(register__n11627) );
  AO22x1_ASAP7_75t_R register___U4854 ( .A1(register__n7822), .A2(register__net125170), .B1(register__n8505), .B2(register__n436), 
        .Y(register__n11506) );
  AO22x1_ASAP7_75t_R register___U4855 ( .A1(register__n9286), .A2(register__n1226), .B1(register__n10169), .B2(register__n75), 
        .Y(register__n10694) );
  AO22x1_ASAP7_75t_R register___U4856 ( .A1(register__net110126), .A2(register__n768), .B1(register__net93440), .B2(
        C6422_net60437), .Y(register__n11010) );
  AO22x1_ASAP7_75t_R register___U4857 ( .A1(register__net112285), .A2(register__n77), .B1(register__net93404), .B2(register__n75), 
        .Y(register__n10713) );
  AO22x1_ASAP7_75t_R register___U4858 ( .A1(register__n6655), .A2(register__n77), .B1(register__n10261), .B2(register__n75), .Y(
        n10991) );
  AO22x1_ASAP7_75t_R register___U4859 ( .A1(register__n6965), .A2(register__n77), .B1(register__n10289), .B2(register__n75), .Y(
        n11031) );
  AO22x1_ASAP7_75t_R register___U4860 ( .A1(register__n9297), .A2(register__n77), .B1(register__n10187), .B2(register__n75), .Y(
        n10652) );
  AO22x1_ASAP7_75t_R register___U4861 ( .A1(register__n9804), .A2(register__net121619), .B1(register__n10203), .B2(
        C6422_net70534), .Y(register__n11119) );
  AO22x1_ASAP7_75t_R register___U4862 ( .A1(register__n10432), .A2(register__net125170), .B1(register__n10428), .B2(
        C6423_net68914), .Y(register__n11355) );
  HB1xp67_ASAP7_75t_R register___U4863 ( .A(register__n11492), .Y(register__n2837) );
  BUFx12f_ASAP7_75t_R register___U4864 ( .A(register__n9366), .Y(register__n9365) );
  INVx1_ASAP7_75t_R register___U4865 ( .A(register__n11249), .Y(register__n1516) );
  INVx1_ASAP7_75t_R register___U4866 ( .A(register__n2078), .Y(register__n1517) );
  INVxp33_ASAP7_75t_R register___U4867 ( .A(register__n2285), .Y(register__n1518) );
  INVx1_ASAP7_75t_R register___U4868 ( .A(register__n1962), .Y(register__n1519) );
  INVx2_ASAP7_75t_R register___U4869 ( .A(register__n1961), .Y(register__n1520) );
  INVxp67_ASAP7_75t_R register___U4870 ( .A(register__n11906), .Y(register__n1521) );
  INVxp33_ASAP7_75t_R register___U4871 ( .A(register__n2286), .Y(register__n1522) );
  INVx1_ASAP7_75t_R register___U4872 ( .A(register__n7088), .Y(register__n1523) );
  INVxp33_ASAP7_75t_R register___U4873 ( .A(register__n11908), .Y(register__n1528) );
  INVx1_ASAP7_75t_R register___U4874 ( .A(register__n1982), .Y(register__n1530) );
  INVx1_ASAP7_75t_R register___U4875 ( .A(register__n1980), .Y(register__n1531) );
  INVx1_ASAP7_75t_R register___U4876 ( .A(register__n1983), .Y(register__n1532) );
  INVx1_ASAP7_75t_R register___U4877 ( .A(register__n11907), .Y(register__n1533) );
  INVx1_ASAP7_75t_R register___U4878 ( .A(register__n2923), .Y(register__n1534) );
  INVx1_ASAP7_75t_R register___U4879 ( .A(register__n2007), .Y(register__n1536) );
  INVx1_ASAP7_75t_R register___U4880 ( .A(register__n2006), .Y(register__n1537) );
  INVx1_ASAP7_75t_R register___U4881 ( .A(register__n2009), .Y(register__n1538) );
  INVx1_ASAP7_75t_R register___U4882 ( .A(register__n2008), .Y(register__n1539) );
  INVx2_ASAP7_75t_R register___U4883 ( .A(register__n11828), .Y(register__n1541) );
  INVx2_ASAP7_75t_R register___U4884 ( .A(register__n6463), .Y(register__n1542) );
  INVx1_ASAP7_75t_R register___U4885 ( .A(register__n6464), .Y(register__n1543) );
  INVx3_ASAP7_75t_R register___U4886 ( .A(register__n4037), .Y(register__n1546) );
  HB1xp67_ASAP7_75t_R register___U4887 ( .A(register__n3716), .Y(register__n4271) );
  CKINVDCx5p33_ASAP7_75t_R register___U4888 ( .A(register__n11907), .Y(register__n1970) );
  BUFx3_ASAP7_75t_R register___U4889 ( .A(register__n2078), .Y(register__n1962) );
  INVx4_ASAP7_75t_R register___U4890 ( .A(register__n1960), .Y(register__n1961) );
  INVxp67_ASAP7_75t_R register___U4891 ( .A(register__n11827), .Y(register__n11906) );
  BUFx6f_ASAP7_75t_R register___U4892 ( .A(register__n7088), .Y(register__n7087) );
  HB1xp67_ASAP7_75t_R register___U4893 ( .A(register__n11908), .Y(register__n2923) );
  INVx2_ASAP7_75t_R register___U4894 ( .A(register__n2005), .Y(register__n2008) );
  INVx6_ASAP7_75t_R register___U4895 ( .A(register__n1970), .Y(register__n1971) );
  BUFx6f_ASAP7_75t_R register___U4896 ( .A(register__n11829), .Y(register__n11828) );
  BUFx6f_ASAP7_75t_R register___U4897 ( .A(register__n11829), .Y(register__n6463) );
  BUFx6f_ASAP7_75t_R register___U4898 ( .A(register__n11829), .Y(register__n6464) );
  BUFx6f_ASAP7_75t_R register___U4899 ( .A(register__n6463), .Y(register__n3159) );
  BUFx6f_ASAP7_75t_R register___U4900 ( .A(register__n11828), .Y(register__n3120) );
  HB1xp67_ASAP7_75t_R register___U4901 ( .A(register__n13233), .Y(register__n3551) );
  HB1xp67_ASAP7_75t_R register___U4902 ( .A(register__n5277), .Y(register__n5276) );
  HB1xp67_ASAP7_75t_R register___U4903 ( .A(register__n10676), .Y(register__n5277) );
  AO22x1_ASAP7_75t_R register___U4904 ( .A1(register__n8815), .A2(register__net125170), .B1(register__n7222), .B2(register__n515), 
        .Y(register__n11647) );
  INVx1_ASAP7_75t_R register___U4905 ( .A(register__n11354), .Y(register__n1555) );
  INVxp67_ASAP7_75t_R register___U4906 ( .A(register__n4393), .Y(register__n4852) );
  HB1xp67_ASAP7_75t_R register___U4907 ( .A(register__n11911), .Y(register__n3716) );
  OA22x2_ASAP7_75t_R register___U4908 ( .A1(register__n1557), .A2(register__n1558), .B1(register__n1559), .B2(register__n1509), 
        .Y(register__n1556) );
  CKINVDCx20_ASAP7_75t_R register___U4909 ( .A(register__n10205), .Y(register__n1559) );
  INVx1_ASAP7_75t_R register___U4910 ( .A(register__n12597), .Y(register__n1560) );
  AO22x1_ASAP7_75t_R register___U4911 ( .A1(register__n9638), .A2(register__net125170), .B1(register__n9949), .B2(
        net94400), .Y(register__n11229) );
  AO22x1_ASAP7_75t_R register___U4912 ( .A1(register__n4958), .A2(register__net125170), .B1(register__n6323), .B2(register__n515), 
        .Y(register__n11208) );
  HB1xp67_ASAP7_75t_R register___U4913 ( .A(register__n11258), .Y(register__n2930) );
  AO22x1_ASAP7_75t_R register___U4914 ( .A1(register__n9589), .A2(register__net93569), .B1(register__n10010), .B2(
        net147378), .Y(register__n11258) );
  HB1xp67_ASAP7_75t_R register___U4915 ( .A(register__n5049), .Y(register__n4376) );
  HB1xp67_ASAP7_75t_R register___U4916 ( .A(register__n5049), .Y(register__n4375) );
  HB1xp67_ASAP7_75t_R register___U4917 ( .A(register__n5531), .Y(register__n11757) );
  BUFx6f_ASAP7_75t_R register___U4918 ( .A(register__n3822), .Y(register__n7663) );
  HB1xp67_ASAP7_75t_R register___U4919 ( .A(register__n11758), .Y(register__n3257) );
  HB1xp67_ASAP7_75t_R register___U4920 ( .A(register__n11760), .Y(register__n11756) );
  HB1xp67_ASAP7_75t_R register___U4921 ( .A(register__n3511), .Y(register__n3509) );
  INVx2_ASAP7_75t_R register___U4922 ( .A(register__n4359), .Y(register__n5702) );
  AO22x1_ASAP7_75t_R register___U4923 ( .A1(register__n10519), .A2(register__net93569), .B1(register__n5207), .B2(
        net147378), .Y(register__n11492) );
  NOR2xp67_ASAP7_75t_R register___U4924 ( .A(register__n519), .B(register__n2458), .Y(register__n2459) );
  BUFx3_ASAP7_75t_R register___U4925 ( .A(register__n1194), .Y(register__n1563) );
  INVxp67_ASAP7_75t_R register___U4926 ( .A(register__net67384), .Y(register__n2149) );
  INVxp67_ASAP7_75t_R register___U4927 ( .A(register__n2142), .Y(register__n2140) );
  CKINVDCx10_ASAP7_75t_R register___U4928 ( .A(register__net67412), .Y(register__net74029) );
  INVx1_ASAP7_75t_R register___U4929 ( .A(register__net73977), .Y(register__net67384) );
  INVxp33_ASAP7_75t_R register___U4930 ( .A(register__n2143), .Y(register__n2144) );
  INVx1_ASAP7_75t_R register___U4931 ( .A(register__n2151), .Y(register__n2152) );
  INVx2_ASAP7_75t_R register___U4932 ( .A(register__net73985), .Y(register__net67382) );
  INVxp67_ASAP7_75t_R register___U4933 ( .A(register__n2149), .Y(register__n2150) );
  INVx1_ASAP7_75t_R register___U4934 ( .A(register__n2147), .Y(register__n2148) );
  BUFx2_ASAP7_75t_R register___U4935 ( .A(register__n4998), .Y(register__n4997) );
  AO22x1_ASAP7_75t_R register___U4936 ( .A1(register__n8761), .A2(register__net125170), .B1(register__n9947), .B2(
        net94399), .Y(register__n11249) );
  BUFx2_ASAP7_75t_R register___U4937 ( .A(register__n6805), .Y(register__n6804) );
  HB1xp67_ASAP7_75t_R register___U4938 ( .A(register__n3717), .Y(register__n11911) );
  HB1xp67_ASAP7_75t_R register___U4939 ( .A(register__n4912), .Y(register__n4911) );
  AO22x1_ASAP7_75t_R register___U4940 ( .A1(register__n9345), .A2(register__net136978), .B1(register__n5835), .B2(
        net138612), .Y(register__n11666) );
  AO22x1_ASAP7_75t_R register___U4941 ( .A1(register__net90793), .A2(register__C6423_net61340), .B1(register__net90041), 
        .B2(register__n334), .Y(register__n11290) );
  AO22x1_ASAP7_75t_R register___U4942 ( .A1(register__n9762), .A2(register__C6423_net61340), .B1(register__n10155), 
        .B2(register__n334), .Y(register__n11313) );
  AOI21xp33_ASAP7_75t_R register___U4943 ( .A1(register__net94399), .A2(register__net88628), .B(register__n1897), .Y(
        n2726) );
  AO22x1_ASAP7_75t_R register___U4944 ( .A1(register__n9911), .A2(register__net125170), .B1(register__n10214), .B2(register__n515), .Y(register__n11417) );
  HB1xp67_ASAP7_75t_R register___U4945 ( .A(register__n12911), .Y(register__n3126) );
  INVx1_ASAP7_75t_R register___U4946 ( .A(register__n11651), .Y(register__n1571) );
  HB1xp67_ASAP7_75t_R register___U4947 ( .A(register__n4587), .Y(register__n1572) );
  INVx1_ASAP7_75t_R register___U4948 ( .A(register__n12866), .Y(register__n1573) );
  INVx1_ASAP7_75t_R register___U4949 ( .A(register__n11885), .Y(register__n4587) );
  INVx1_ASAP7_75t_R register___U4950 ( .A(register__n2815), .Y(register__n1945) );
  INVx1_ASAP7_75t_R register___U4951 ( .A(register__n2812), .Y(register__n1933) );
  INVx1_ASAP7_75t_R register___U4952 ( .A(register__n2810), .Y(register__n1926) );
  INVx1_ASAP7_75t_R register___U4953 ( .A(register__n2805), .Y(register__n1952) );
  INVx1_ASAP7_75t_R register___U4954 ( .A(register__n2805), .Y(register__n2816) );
  INVx2_ASAP7_75t_R register___U4955 ( .A(register__n1968), .Y(register__n2809) );
  INVxp33_ASAP7_75t_R register___U4956 ( .A(register__n12498), .Y(register__n2983) );
  BUFx2_ASAP7_75t_R register___U4957 ( .A(register__n2804), .Y(register__n2813) );
  INVx1_ASAP7_75t_R register___U4958 ( .A(register__n1930), .Y(register__n1927) );
  INVx1_ASAP7_75t_R register___U4959 ( .A(register__n1945), .Y(register__n1942) );
  INVx1_ASAP7_75t_R register___U4960 ( .A(register__n1941), .Y(register__n1938) );
  INVx1_ASAP7_75t_R register___U4961 ( .A(register__n1933), .Y(register__n1931) );
  INVx1_ASAP7_75t_R register___U4962 ( .A(register__n1926), .Y(register__n1923) );
  BUFx2_ASAP7_75t_R register___U4963 ( .A(register__n2802), .Y(register__n1968) );
  INVx1_ASAP7_75t_R register___U4964 ( .A(register__n2809), .Y(register__n1921) );
  INVx1_ASAP7_75t_R register___U4965 ( .A(register__n2816), .Y(register__n2819) );
  INVxp67_ASAP7_75t_R register___U4966 ( .A(register__n2817), .Y(register__n2806) );
  INVx1_ASAP7_75t_R register___U4967 ( .A(register__n1952), .Y(register__n1957) );
  HB1xp67_ASAP7_75t_R register___U4968 ( .A(register__n9408), .Y(register__n5734) );
  HB1xp67_ASAP7_75t_R register___U4969 ( .A(register__n11590), .Y(register__n6805) );
  AO22x1_ASAP7_75t_R register___U4970 ( .A1(register__n9834), .A2(register__C6423_net61318), .B1(register__n6644), .B2(
        n1447), .Y(register__n11590) );
  OAI22xp33_ASAP7_75t_R register___U4971 ( .A1(register__net62826), .A2(register__n1568), .B1(register__net88760), .B2(
        n1193), .Y(register__n1574) );
  INVxp33_ASAP7_75t_R register___U4972 ( .A(register__n4271), .Y(register__n11908) );
  HB1xp67_ASAP7_75t_R register___U4973 ( .A(register__n12599), .Y(register__n3858) );
  INVx2_ASAP7_75t_R register___U4974 ( .A(register__net62866), .Y(register__net62832) );
  HB1xp67_ASAP7_75t_R register___U4975 ( .A(register__n4394), .Y(register__n4393) );
  HB1xp67_ASAP7_75t_R register___U4976 ( .A(register__n11667), .Y(register__n4912) );
  HB1xp67_ASAP7_75t_R register___U4977 ( .A(register__net64732), .Y(register__net64696) );
  HB1xp67_ASAP7_75t_R register___U4978 ( .A(register__n12571), .Y(register__n4418) );
  AO22x1_ASAP7_75t_R register___U4979 ( .A1(register__n9266), .A2(register__C6423_net68948), .B1(register__n10319), 
        .B2(register__net120961), .Y(register__n11460) );
  HB1xp67_ASAP7_75t_R register___U4980 ( .A(register__n11449), .Y(register__n7016) );
  HB1xp67_ASAP7_75t_R register___U4981 ( .A(register__n13002), .Y(register__n4083) );
  HB1xp67_ASAP7_75t_R register___U4982 ( .A(register__n11049), .Y(register__n4998) );
  AO22x1_ASAP7_75t_R register___U4983 ( .A1(register__n9296), .A2(register__n933), .B1(register__n10446), .B2(register__n1906), 
        .Y(register__n11193) );
  AO22x1_ASAP7_75t_R register___U4984 ( .A1(register__n8781), .A2(register__net126316), .B1(register__net123880), .B2(
        n10325), .Y(register__n11137) );
  INVxp67_ASAP7_75t_R register___U4985 ( .A(register__n5572), .Y(register__n8658) );
  HB1xp67_ASAP7_75t_R register___U4986 ( .A(register__n5573), .Y(register__n5572) );
  HB1xp67_ASAP7_75t_R register___U4987 ( .A(register__n12530), .Y(register__n5776) );
  HB1xp67_ASAP7_75t_R register___U4988 ( .A(register__n12601), .Y(register__n4394) );
  AO22x1_ASAP7_75t_R register___U4989 ( .A1(register__n7540), .A2(register__net131160), .B1(register__n10323), .B2(
        net120912), .Y(register__n11049) );
  HB1xp67_ASAP7_75t_R register___U4990 ( .A(register__n12877), .Y(register__n5573) );
  HB1xp67_ASAP7_75t_R register___U4991 ( .A(register__n7353), .Y(register__n7352) );
  HB1xp67_ASAP7_75t_R register___U4992 ( .A(register__n12972), .Y(register__n2949) );
  AND2x2_ASAP7_75t_R register___U4993 ( .A(register__n7595), .B(register__n7594), .Y(register__n1582) );
  INVx2_ASAP7_75t_R register___U4994 ( .A(register__n11404), .Y(register__n3792) );
  HB1xp67_ASAP7_75t_R register___U4995 ( .A(register__n12740), .Y(register__n3772) );
  INVx1_ASAP7_75t_R register___U4996 ( .A(register__n10909), .Y(register__n8697) );
  BUFx3_ASAP7_75t_R register___U4997 ( .A(register__n11506), .Y(register__n4028) );
  AO22x1_ASAP7_75t_R register___U4998 ( .A1(register__n9579), .A2(register__n309), .B1(register__n9999), .B2(
        C6423_net74857), .Y(register__n11578) );
  INVx1_ASAP7_75t_R register___U4999 ( .A(register__n10779), .Y(register__n2254) );
  INVxp67_ASAP7_75t_R register___U5000 ( .A(register__n13065), .Y(register__n8685) );
  INVxp67_ASAP7_75t_R register___U5001 ( .A(register__n3022), .Y(register__n1585) );
  INVxp67_ASAP7_75t_R register___U5002 ( .A(register__n3071), .Y(register__n1587) );
  INVxp67_ASAP7_75t_R register___U5003 ( .A(register__n3071), .Y(register__n1588) );
  INVxp33_ASAP7_75t_R register___U5004 ( .A(register__n3071), .Y(register__n1592) );
  INVx1_ASAP7_75t_R register___U5005 ( .A(register__n2935), .Y(register__n1597) );
  INVx2_ASAP7_75t_R register___U5006 ( .A(register__n2935), .Y(register__n1600) );
  INVx1_ASAP7_75t_R register___U5007 ( .A(register__n11895), .Y(register__n1601) );
  INVx2_ASAP7_75t_R register___U5008 ( .A(register__n11817), .Y(register__n1605) );
  INVx2_ASAP7_75t_R register___U5009 ( .A(register__n3072), .Y(register__n11895) );
  HB1xp67_ASAP7_75t_R register___U5010 ( .A(register__n12850), .Y(register__n6790) );
  HB1xp67_ASAP7_75t_R register___U5011 ( .A(register__n12846), .Y(register__n4878) );
  HB1xp67_ASAP7_75t_R register___U5012 ( .A(register__n12841), .Y(register__n5005) );
  HB1xp67_ASAP7_75t_R register___U5013 ( .A(register__n12833), .Y(register__n5098) );
  HB1xp67_ASAP7_75t_R register___U5014 ( .A(register__n4414), .Y(register__n4413) );
  HB1xp67_ASAP7_75t_R register___U5015 ( .A(register__n13179), .Y(register__n4414) );
  BUFx6f_ASAP7_75t_R register___U5016 ( .A(register__net140665), .Y(register__net140664) );
  AND3x1_ASAP7_75t_R register___U5017 ( .A(register__n7272), .B(register__n7271), .C(register__n7875), .Y(register__n2798) );
  HB1xp67_ASAP7_75t_R register___U5018 ( .A(register__n12720), .Y(register__n4542) );
  HB1xp67_ASAP7_75t_R register___U5019 ( .A(register__n3842), .Y(register__n5223) );
  AO22x1_ASAP7_75t_R register___U5020 ( .A1(register__n5192), .A2(register__net93569), .B1(register__n10003), .B2(
        C6423_net74857), .Y(register__n11538) );
  OAI22xp5_ASAP7_75t_R register___U5021 ( .A1(register__n53), .A2(register__n7889), .B1(register__net61369), .B2(
        net62848), .Y(read_reg_data_1[29]) );
  HB1xp67_ASAP7_75t_R register___U5022 ( .A(register__n12860), .Y(register__n4077) );
  HB1xp67_ASAP7_75t_R register___U5023 ( .A(register__n4784), .Y(register__n4783) );
  HB1xp67_ASAP7_75t_R register___U5024 ( .A(register__n12926), .Y(register__n4784) );
  AO22x1_ASAP7_75t_R register___U5025 ( .A1(register__n9754), .A2(register__net93569), .B1(register__n10148), .B2(
        C6423_net74857), .Y(register__n11404) );
  INVx4_ASAP7_75t_R register___U5026 ( .A(register__n11306), .Y(register__n9148) );
  INVx2_ASAP7_75t_R register___U5027 ( .A(register__n1968), .Y(register__n2808) );
  AO22x1_ASAP7_75t_R register___U5028 ( .A1(register__n9597), .A2(register__n128), .B1(register__n10018), .B2(register__n1444), 
        .Y(register__n11570) );
  AOI22xp33_ASAP7_75t_R register___U5029 ( .A1(register__net130838), .A2(register__n1943), .B1(register__C6422_net59961), .B2(register__n2814), .Y(register__n12874) );
  INVx1_ASAP7_75t_R register___U5030 ( .A(register__n2811), .Y(register__n1930) );
  INVx1_ASAP7_75t_R register___U5031 ( .A(register__n12861), .Y(register__n1609) );
  HB1xp67_ASAP7_75t_R register___U5032 ( .A(register__n12864), .Y(register__n3397) );
  INVx1_ASAP7_75t_R register___U5033 ( .A(register__n11438), .Y(register__n1610) );
  HB1xp67_ASAP7_75t_R register___U5034 ( .A(register__n3842), .Y(register__n12478) );
  INVxp33_ASAP7_75t_R register___U5035 ( .A(register__n12498), .Y(register__n2802) );
  AOI22xp33_ASAP7_75t_R register___U5036 ( .A1(register__n6925), .A2(register__n1867), .B1(register__n6375), .B2(register__n1348), 
        .Y(register__n1611) );
  INVx6_ASAP7_75t_R register___U5037 ( .A(register__n3730), .Y(register__n12433) );
  AO22x1_ASAP7_75t_R register___U5038 ( .A1(register__n5191), .A2(register__n1771), .B1(register__n10003), .B2(
        net126625), .Y(register__n10927) );
  INVx2_ASAP7_75t_R register___U5039 ( .A(register__n11112), .Y(register__n6457) );
  HB1xp67_ASAP7_75t_R register___U5040 ( .A(register__n284), .Y(register__C6423_net74851) );
  AO22x1_ASAP7_75t_R register___U5041 ( .A1(register__n7437), .A2(register__net125170), .B1(register__n6562), .B2(register__n515), 
        .Y(register__n11484) );
  BUFx3_ASAP7_75t_R register___U5042 ( .A(register__n3256), .Y(register__n3189) );
  HB1xp67_ASAP7_75t_R register___U5043 ( .A(register__n12734), .Y(register__n3461) );
  INVx1_ASAP7_75t_R register___U5044 ( .A(register__n12881), .Y(register__n1612) );
  HB1xp67_ASAP7_75t_R register___U5045 ( .A(register__n12623), .Y(register__n4668) );
  INVxp67_ASAP7_75t_R register___U5046 ( .A(register__n3930), .Y(register__n6437) );
  HB1xp67_ASAP7_75t_R register___U5047 ( .A(register__n3931), .Y(register__n3930) );
  INVx1_ASAP7_75t_R register___U5048 ( .A(register__n11308), .Y(register__n1613) );
  INVx1_ASAP7_75t_R register___U5049 ( .A(register__n10748), .Y(register__n1614) );
  INVx6_ASAP7_75t_R register___U5050 ( .A(register__n3255), .Y(register__n12143) );
  AO22x1_ASAP7_75t_R register___U5051 ( .A1(register__n9688), .A2(register__C6422_net60422), .B1(register__n9959), .B2(
        net123857), .Y(register__n10876) );
  AOI22xp33_ASAP7_75t_R register___U5052 ( .A1(register__n12211), .A2(register__n4579), .B1(register__n1615), .B2(register__n1120), .Y(register__n13075) );
  CKINVDCx20_ASAP7_75t_R register___U5053 ( .A(register__n9335), .Y(register__n1615) );
  INVxp67_ASAP7_75t_R register___U5054 ( .A(register__n3955), .Y(register__n6134) );
  HB1xp67_ASAP7_75t_R register___U5055 ( .A(register__n12936), .Y(register__n3955) );
  INVxp67_ASAP7_75t_R register___U5056 ( .A(register__n1793), .Y(register__n1619) );
  INVxp33_ASAP7_75t_R register___U5057 ( .A(register__n1644), .Y(register__n1623) );
  INVxp67_ASAP7_75t_R register___U5058 ( .A(register__n1776), .Y(register__n1626) );
  INVx2_ASAP7_75t_R register___U5059 ( .A(register__n1778), .Y(register__n1627) );
  INVx1_ASAP7_75t_R register___U5060 ( .A(register__n1782), .Y(register__n1628) );
  INVx1_ASAP7_75t_R register___U5061 ( .A(register__n1780), .Y(register__n1634) );
  INVx1_ASAP7_75t_R register___U5062 ( .A(register__n1786), .Y(register__n1637) );
  INVx2_ASAP7_75t_R register___U5063 ( .A(register__n1789), .Y(register__n1638) );
  INVx2_ASAP7_75t_R register___U5064 ( .A(register__n1791), .Y(register__n1639) );
  INVx2_ASAP7_75t_R register___U5065 ( .A(register__n3043), .Y(register__n1640) );
  INVxp67_ASAP7_75t_R register___U5066 ( .A(register__n11893), .Y(register__n1781) );
  INVx1_ASAP7_75t_R register___U5067 ( .A(register__n11892), .Y(register__n1785) );
  INVxp33_ASAP7_75t_R register___U5068 ( .A(register__n1775), .Y(register__n1776) );
  INVx2_ASAP7_75t_R register___U5069 ( .A(register__n1777), .Y(register__n1778) );
  INVxp67_ASAP7_75t_R register___U5070 ( .A(register__n1781), .Y(register__n1782) );
  INVxp67_ASAP7_75t_R register___U5071 ( .A(register__n1779), .Y(register__n1780) );
  INVx1_ASAP7_75t_R register___U5072 ( .A(register__n11810), .Y(register__n11892) );
  INVx2_ASAP7_75t_R register___U5073 ( .A(register__n1618), .Y(register__n1787) );
  INVx2_ASAP7_75t_R register___U5074 ( .A(register__n1788), .Y(register__n1789) );
  INVx2_ASAP7_75t_R register___U5075 ( .A(register__n1790), .Y(register__n1791) );
  INVx1_ASAP7_75t_R register___U5076 ( .A(register__n12210), .Y(register__n12196) );
  INVx1_ASAP7_75t_R register___U5077 ( .A(register__n12209), .Y(register__n12195) );
  INVxp67_ASAP7_75t_R register___U5078 ( .A(register__n1887), .Y(register__n2826) );
  HB1xp67_ASAP7_75t_R register___U5079 ( .A(register__n12862), .Y(register__n3662) );
  HB1xp67_ASAP7_75t_R register___U5080 ( .A(register__n12884), .Y(register__n5569) );
  HB1xp67_ASAP7_75t_R register___U5081 ( .A(register__n12878), .Y(register__n3933) );
  HB1xp67_ASAP7_75t_R register___U5082 ( .A(register__n12887), .Y(register__n3923) );
  OAI21xp33_ASAP7_75t_R register___U5083 ( .A1(register__net103314), .A2(register__net130087), .B(register__n17), .Y(
        n2661) );
  AO22x1_ASAP7_75t_R register___U5084 ( .A1(register__net109927), .A2(register__net110414), .B1(register__net89413), 
        .B2(register__n1073), .Y(register__n11613) );
  AO22x1_ASAP7_75t_R register___U5085 ( .A1(register__n8813), .A2(register__C6423_net61340), .B1(register__n8821), .B2(
        n334), .Y(register__n11651) );
  INVx1_ASAP7_75t_R register___U5086 ( .A(register__n11025), .Y(register__n1648) );
  INVxp67_ASAP7_75t_R register___U5087 ( .A(register__n12760), .Y(register__n6132) );
  INVxp67_ASAP7_75t_R register___U5088 ( .A(register__n4308), .Y(register__n7924) );
  HB1xp67_ASAP7_75t_R register___U5089 ( .A(register__n4309), .Y(register__n4308) );
  HB1xp67_ASAP7_75t_R register___U5090 ( .A(register__n11550), .Y(register__n4309) );
  AO22x1_ASAP7_75t_R register___U5091 ( .A1(register__n8759), .A2(register__net125169), .B1(register__n9945), .B2(register__n515), 
        .Y(register__n11550) );
  NAND2xp33_ASAP7_75t_R register___U5092 ( .A(register__net89589), .B(register__C6422_net70534), .Y(register__n1841) );
  AO22x1_ASAP7_75t_R register___U5093 ( .A1(register__n9754), .A2(register__net118635), .B1(register__n10148), .B2(
        net126625), .Y(register__n10777) );
  AO22x1_ASAP7_75t_R register___U5094 ( .A1(register__n9857), .A2(register__n387), .B1(register__n10327), .B2(register__net120912), .Y(register__n11139) );
  AND2x2_ASAP7_75t_R register___U5095 ( .A(register__n10860), .B(register__n7884), .Y(register__n1649) );
  AND3x1_ASAP7_75t_R register___U5096 ( .A(register__n1649), .B(register__n764), .C(register__n10861), .Y(register__n4032) );
  INVxp67_ASAP7_75t_R register___U5097 ( .A(register__n13095), .Y(register__n8654) );
  INVx1_ASAP7_75t_R register___U5098 ( .A(register__net110413), .Y(register__n1650) );
  HB1xp67_ASAP7_75t_R register___U5099 ( .A(register__net110413), .Y(register__net110412) );
  HB1xp67_ASAP7_75t_R register___U5100 ( .A(register__n3325), .Y(register__n11742) );
  BUFx12f_ASAP7_75t_R register___U5101 ( .A(register__n3382), .Y(register__n3381) );
  HB1xp67_ASAP7_75t_R register___U5102 ( .A(register__n3380), .Y(register__n5500) );
  BUFx4f_ASAP7_75t_R register___U5103 ( .A(register__n3326), .Y(register__n5640) );
  BUFx6f_ASAP7_75t_R register___U5104 ( .A(register__n5640), .Y(register__n11743) );
  BUFx12f_ASAP7_75t_R register___U5105 ( .A(register__n3879), .Y(register__n3264) );
  BUFx12f_ASAP7_75t_R register___U5106 ( .A(register__n8336), .Y(register__n3823) );
  BUFx12f_ASAP7_75t_R register___U5107 ( .A(register__n3937), .Y(register__n3946) );
  INVx6_ASAP7_75t_R register___U5108 ( .A(register__n4637), .Y(register__n11859) );
  INVx4_ASAP7_75t_R register___U5109 ( .A(register__n3823), .Y(register__n11860) );
  AO22x1_ASAP7_75t_R register___U5110 ( .A1(register__n9603), .A2(register__n40), .B1(register__n9427), .B2(
        C6422_net60399), .Y(register__n10603) );
  INVx6_ASAP7_75t_R register___U5111 ( .A(register__net137417), .Y(register__n1651) );
  AO22x1_ASAP7_75t_R register___U5112 ( .A1(register__n9664), .A2(register__n1867), .B1(register__net96692), .B2(register__n9993), 
        .Y(register__n10624) );
  AO22x1_ASAP7_75t_R register___U5113 ( .A1(register__n9666), .A2(register__net91683), .B1(register__n9425), .B2(
        net96692), .Y(register__n10579) );
  AOI21xp33_ASAP7_75t_R register___U5114 ( .A1(register__C6423_net68950), .A2(register__net93468), .B(register__n2556), 
        .Y(register__n2580) );
  AO22x1_ASAP7_75t_R register___U5115 ( .A1(register__n8797), .A2(register__C6423_net61326), .B1(register__n9131), .B2(
        n2138), .Y(register__n11710) );
  AO22x1_ASAP7_75t_R register___U5116 ( .A1(register__n9268), .A2(register__C6423_net61326), .B1(register__n10191), 
        .B2(register__n1999), .Y(register__n11688) );
  INVx2_ASAP7_75t_R register___U5117 ( .A(register__n4573), .Y(register__n7920) );
  AND4x1_ASAP7_75t_R register___U5118 ( .A(register__n6193), .B(register__n6191), .C(register__n6192), .D(register__n3167), .Y(
        n10908) );
  INVxp67_ASAP7_75t_R register___U5119 ( .A(register__n2120), .Y(register__n1658) );
  INVxp33_ASAP7_75t_R register___U5120 ( .A(register__net66594), .Y(register__n1662) );
  INVx1_ASAP7_75t_R register___U5121 ( .A(register__n2122), .Y(register__n1663) );
  INVxp67_ASAP7_75t_R register___U5122 ( .A(register__n2094), .Y(register__n1665) );
  INVx2_ASAP7_75t_R register___U5123 ( .A(register__n2116), .Y(register__n1666) );
  INVx1_ASAP7_75t_R register___U5124 ( .A(register__n2096), .Y(register__n1667) );
  INVxp33_ASAP7_75t_R register___U5125 ( .A(register__net73061), .Y(register__n1668) );
  INVx1_ASAP7_75t_R register___U5126 ( .A(register__net73059), .Y(register__n1669) );
  INVx1_ASAP7_75t_R register___U5127 ( .A(register__net104558), .Y(register__n1670) );
  INVx1_ASAP7_75t_R register___U5128 ( .A(register__net104559), .Y(register__n1671) );
  INVxp67_ASAP7_75t_R register___U5129 ( .A(register__n2098), .Y(register__n1672) );
  INVx1_ASAP7_75t_R register___U5130 ( .A(register__n2100), .Y(register__n1673) );
  INVx1_ASAP7_75t_R register___U5131 ( .A(register__net66582), .Y(register__n1674) );
  INVx1_ASAP7_75t_R register___U5132 ( .A(register__n2104), .Y(register__n1675) );
  INVx1_ASAP7_75t_R register___U5133 ( .A(register__n2102), .Y(register__n1676) );
  INVx1_ASAP7_75t_R register___U5134 ( .A(register__n2108), .Y(register__n1678) );
  INVx1_ASAP7_75t_R register___U5135 ( .A(register__n2106), .Y(register__n1679) );
  INVx1_ASAP7_75t_R register___U5136 ( .A(register__n2110), .Y(register__n1681) );
  INVx1_ASAP7_75t_R register___U5137 ( .A(register__n2114), .Y(register__n1682) );
  INVx1_ASAP7_75t_R register___U5138 ( .A(register__n2112), .Y(register__n1683) );
  INVxp33_ASAP7_75t_R register___U5139 ( .A(register__net130481), .Y(register__n2120) );
  INVxp33_ASAP7_75t_R register___U5140 ( .A(register__n2093), .Y(register__n2094) );
  INVx1_ASAP7_75t_R register___U5141 ( .A(register__n2095), .Y(register__n2096) );
  BUFx6f_ASAP7_75t_R register___U5142 ( .A(register__net73061), .Y(register__net104558) );
  INVxp33_ASAP7_75t_R register___U5143 ( .A(register__n2097), .Y(register__n2098) );
  INVx1_ASAP7_75t_R register___U5144 ( .A(register__n2099), .Y(register__n2100) );
  INVx1_ASAP7_75t_R register___U5145 ( .A(register__n2101), .Y(register__n2102) );
  BUFx12f_ASAP7_75t_R register___U5146 ( .A(register__net104559), .Y(register__net137800) );
  INVx1_ASAP7_75t_R register___U5147 ( .A(register__n2111), .Y(register__n2112) );
  INVx3_ASAP7_75t_R register___U5148 ( .A(register__n2122), .Y(register__n2115) );
  INVxp67_ASAP7_75t_R register___U5149 ( .A(register__net146710), .Y(register__n2095) );
  INVx1_ASAP7_75t_R register___U5150 ( .A(register__net73059), .Y(register__n2099) );
  INVx1_ASAP7_75t_R register___U5151 ( .A(register__net104559), .Y(register__n2101) );
  INVx1_ASAP7_75t_R register___U5152 ( .A(register__net66582), .Y(register__n2107) );
  INVx2_ASAP7_75t_R register___U5153 ( .A(register__net137800), .Y(register__n2109) );
  INVx4_ASAP7_75t_R register___U5154 ( .A(register__net137800), .Y(register__net73019) );
  INVx1_ASAP7_75t_R register___U5155 ( .A(register__net66574), .Y(register__n2113) );
  INVx1_ASAP7_75t_R register___U5156 ( .A(register__n11270), .Y(register__n1685) );
  INVxp67_ASAP7_75t_R register___U5157 ( .A(register__n4462), .Y(register__n6151) );
  HB1xp67_ASAP7_75t_R register___U5158 ( .A(register__n4463), .Y(register__n4462) );
  HB1xp67_ASAP7_75t_R register___U5159 ( .A(register__n4227), .Y(register__n4226) );
  INVxp67_ASAP7_75t_R register___U5160 ( .A(register__n4226), .Y(register__n6747) );
  HB1xp67_ASAP7_75t_R register___U5161 ( .A(register__net147379), .Y(register__C6423_net74855) );
  AO22x1_ASAP7_75t_R register___U5162 ( .A1(register__n9768), .A2(register__net129747), .B1(register__n10110), .B2(
        net139537), .Y(register__n10748) );
  BUFx12f_ASAP7_75t_R register___U5163 ( .A(register__n4848), .Y(register__n3393) );
  INVx6_ASAP7_75t_R register___U5164 ( .A(register__n3393), .Y(register__n12152) );
  HB1xp67_ASAP7_75t_R register___U5165 ( .A(register__n11440), .Y(register__n4227) );
  AO22x1_ASAP7_75t_R register___U5166 ( .A1(register__n8781), .A2(register__C6423_net61343), .B1(register__n10325), 
        .B2(register__net129787), .Y(register__n11715) );
  INVxp67_ASAP7_75t_R register___U5167 ( .A(register__n3037), .Y(register__n6193) );
  HB1xp67_ASAP7_75t_R register___U5168 ( .A(register__n3038), .Y(register__n3037) );
  HB1xp67_ASAP7_75t_R register___U5169 ( .A(register__n10919), .Y(register__n3038) );
  OAI22xp33_ASAP7_75t_R register___U5170 ( .A1(register__net64834), .A2(register__n11860), .B1(register__net89813), 
        .B2(register__n3325), .Y(register__n1686) );
  AOI21xp33_ASAP7_75t_R register___U5171 ( .A1(register__net110412), .A2(register__net90225), .B(register__n2573), .Y(
        n2575) );
  HB1xp67_ASAP7_75t_R register___U5172 ( .A(register__n11316), .Y(register__n4463) );
  AND4x1_ASAP7_75t_R register___U5173 ( .A(register__n5521), .B(register__n5522), .C(register__n8037), .D(register__n4244), .Y(
        n10716) );
  INVx2_ASAP7_75t_R register___U5174 ( .A(register__n3141), .Y(register__n5230) );
  AO22x1_ASAP7_75t_R register___U5175 ( .A1(register__n7520), .A2(register__net91683), .B1(register__n10136), .B2(register__n1356), .Y(register__n11069) );
  HB1xp67_ASAP7_75t_R register___U5176 ( .A(register__n10874), .Y(register__n3093) );
  BUFx6f_ASAP7_75t_R register___U5177 ( .A(register__net66618), .Y(register__net130481) );
  AO22x1_ASAP7_75t_R register___U5178 ( .A1(register__n9110), .A2(register__net91683), .B1(register__n10283), .B2(register__n1359), .Y(register__n11025) );
  INVxp67_ASAP7_75t_R register___U5179 ( .A(register__n4659), .Y(register__n6436) );
  HB1xp67_ASAP7_75t_R register___U5180 ( .A(register__n4660), .Y(register__n4659) );
  BUFx4f_ASAP7_75t_R register___U5181 ( .A(register__net102299), .Y(register__net102304) );
  INVx4_ASAP7_75t_R register___U5182 ( .A(register__net102304), .Y(register__n_cell_124938_net165675) );
  INVx1_ASAP7_75t_R register___U5183 ( .A(register__n13304), .Y(register__n1689) );
  AO22x1_ASAP7_75t_R register___U5184 ( .A1(register__n9724), .A2(register__net129017), .B1(register__n10175), .B2(register__n422), .Y(register__n11466) );
  AO22x1_ASAP7_75t_R register___U5185 ( .A1(register__net90877), .A2(register__n1867), .B1(register__net89969), .B2(
        n1353), .Y(register__n11004) );
  NAND2xp33_ASAP7_75t_R register___U5186 ( .A(register__n1344), .B(register__net89425), .Y(register__n2667) );
  AOI22xp5_ASAP7_75t_R register___U5187 ( .A1(register__n12298), .A2(register__register__n1186), .B1(register__n1690), .B2(register__n118), 
        .Y(register__n13096) );
  CKINVDCx20_ASAP7_75t_R register___U5188 ( .A(register__n8831), .Y(register__n1690) );
  INVx2_ASAP7_75t_R register___U5189 ( .A(register__n12298), .Y(register__n12284) );
  INVxp67_ASAP7_75t_R register___U5190 ( .A(register__n12639), .Y(register__n7085) );
  INVxp33_ASAP7_75t_R register___U5191 ( .A(register__n1836), .Y(register__n1693) );
  INVxp33_ASAP7_75t_R register___U5192 ( .A(register__n1836), .Y(register__n1697) );
  INVxp33_ASAP7_75t_R register___U5193 ( .A(register__n1693), .Y(register__n1708) );
  INVx1_ASAP7_75t_R register___U5194 ( .A(register__n1714), .Y(register__n1715) );
  BUFx12f_ASAP7_75t_R register___U5195 ( .A(register__n6160), .Y(register__n11871) );
  AO22x1_ASAP7_75t_R register___U5196 ( .A1(register__n10481), .A2(register__C6423_net61343), .B1(register__n10462), 
        .B2(register__net122313), .Y(register__n11440) );
  BUFx3_ASAP7_75t_R register___U5197 ( .A(register__n10784), .Y(register__n5473) );
  AO22x1_ASAP7_75t_R register___U5198 ( .A1(register__n9686), .A2(register__C6423_net61340), .B1(register__n9957), .B2(
        net125365), .Y(register__n11533) );
  HB1xp67_ASAP7_75t_R register___U5199 ( .A(register__n11593), .Y(register__n4717) );
  AO22x1_ASAP7_75t_R register___U5200 ( .A1(register__n9682), .A2(register__C6423_net61340), .B1(register__n9953), .B2(
        n334), .Y(register__n11573) );
  AO22x1_ASAP7_75t_R register___U5201 ( .A1(register__n9718), .A2(register__C6423_net61340), .B1(register__n10094), 
        .B2(register__net125365), .Y(register__n11399) );
  INVxp67_ASAP7_75t_R register___U5202 ( .A(register__n11592), .Y(register__n6713) );
  AO22x1_ASAP7_75t_R register___U5203 ( .A1(register__n9714), .A2(register__net131160), .B1(register__n10044), .B2(
        net120912), .Y(register__n10627) );
  INVx2_ASAP7_75t_R register___U5204 ( .A(register__n10737), .Y(register__n8318) );
  AO22x1_ASAP7_75t_R register___U5205 ( .A1(register__n9716), .A2(register__n387), .B1(register__n10046), .B2(register__net120912), .Y(register__n10607) );
  AO22x1_ASAP7_75t_R register___U5206 ( .A1(register__n9778), .A2(register__net110414), .B1(register__n10164), .B2(
        n1074), .Y(register__n11316) );
  AO22x1_ASAP7_75t_R register___U5207 ( .A1(register__n8775), .A2(register__net110414), .B1(register__n10144), .B2(
        n1073), .Y(register__n11382) );
  INVx2_ASAP7_75t_R register___U5208 ( .A(register__n5472), .Y(register__n9226) );
  AOI222xp33_ASAP7_75t_R register___U5209 ( .A1(register__C6422_net59546), .A2(register__n1740), .B1(
        C6422_net59548), .B2(register__n10916), .C1(register__n1580), .C2(register__n9471), .Y(register__n10910) );
  INVx2_ASAP7_75t_R register___U5210 ( .A(register__n10916), .Y(register__n9157) );
  INVx1_ASAP7_75t_R register___U5211 ( .A(register__n9471), .Y(register__n11527) );
  AO22x1_ASAP7_75t_R register___U5212 ( .A1(register__n9613), .A2(register__net126316), .B1(register__n10080), .B2(
        net123880), .Y(register__n10875) );
  AO22x1_ASAP7_75t_R register___U5213 ( .A1(register__n9824), .A2(register__n387), .B1(register__n10235), .B2(register__net120912), .Y(register__n10900) );
  AO22x1_ASAP7_75t_R register___U5214 ( .A1(register__n8929), .A2(register__n387), .B1(register__n10038), .B2(register__net120912), .Y(register__n10877) );
  AO22x1_ASAP7_75t_R register___U5215 ( .A1(register__n8161), .A2(register__net126316), .B1(register__n10158), .B2(
        net123880), .Y(register__n10898) );
  AO22x1_ASAP7_75t_R register___U5216 ( .A1(register__n9770), .A2(register__net126316), .B1(register__n10120), .B2(
        net123880), .Y(register__n10851) );
  AO22x1_ASAP7_75t_R register___U5217 ( .A1(register__n9760), .A2(register__net91683), .B1(register__n10245), .B2(register__n90), 
        .Y(register__n10897) );
  HB1xp67_ASAP7_75t_R register___U5218 ( .A(register__n10670), .Y(register__n4104) );
  AO22x1_ASAP7_75t_R register___U5219 ( .A1(register__n10483), .A2(register__net126316), .B1(register__n10463), .B2(
        net123880), .Y(register__n10670) );
  AO22x1_ASAP7_75t_R register___U5220 ( .A1(register__n9684), .A2(register__C6423_net61340), .B1(register__n9955), .B2(
        n334), .Y(register__n11554) );
  INVx1_ASAP7_75t_R register___U5221 ( .A(register__n10796), .Y(register__n1741) );
  AO22x1_ASAP7_75t_R register___U5222 ( .A1(register__n9262), .A2(register__net126316), .B1(register__n10102), .B2(
        net123880), .Y(register__n10771) );
  NOR2xp67_ASAP7_75t_R register___U5223 ( .A(register__n1687), .B(register__net62848), .Y(register__n2558) );
  AO22x1_ASAP7_75t_R register___U5224 ( .A1(register__net90997), .A2(register__net122249), .B1(register__net89713), 
        .B2(register__net122313), .Y(register__n11270) );
  NOR2xp67_ASAP7_75t_R register___U5225 ( .A(register__n1687), .B(register__net64360), .Y(register__n2614) );
  AO22x1_ASAP7_75t_R register___U5226 ( .A1(register__n9843), .A2(register__C6423_net61340), .B1(register__n10122), 
        .B2(register__net125365), .Y(register__n11593) );
  INVxp67_ASAP7_75t_R register___U5227 ( .A(register__n4389), .Y(register__n6057) );
  HB1xp67_ASAP7_75t_R register___U5228 ( .A(register__n4390), .Y(register__n4389) );
  AO22x1_ASAP7_75t_R register___U5229 ( .A1(register__n9244), .A2(register__net122579), .B1(register__n10444), .B2(
        n1998), .Y(register__n11237) );
  NAND2xp5_ASAP7_75t_R register___U5230 ( .A(register__n1743), .B(register__n1742), .Y(register__n13388) );
  OR2x2_ASAP7_75t_R register___U5231 ( .A(register__n2134), .B(register__n49), .Y(register__n1743) );
  AO22x1_ASAP7_75t_R register___U5232 ( .A1(register__net90713), .A2(register__net126316), .B1(register__net89657), 
        .B2(register__net123880), .Y(register__n10725) );
  INVx2_ASAP7_75t_R register___U5233 ( .A(register__n4245), .Y(register__n5521) );
  HB1xp67_ASAP7_75t_R register___U5234 ( .A(register__n3185), .Y(register__n11772) );
  HB1xp67_ASAP7_75t_R register___U5235 ( .A(register__n3248), .Y(register__n11774) );
  HB1xp67_ASAP7_75t_R register___U5236 ( .A(register__n11771), .Y(register__n11773) );
  HB1xp67_ASAP7_75t_R register___U5237 ( .A(register__n11780), .Y(register__n11775) );
  INVxp67_ASAP7_75t_R register___U5238 ( .A(register__n2012), .Y(register__n1919) );
  HB1xp67_ASAP7_75t_R register___U5239 ( .A(register__n11769), .Y(register__n11770) );
  HB1xp67_ASAP7_75t_R register___U5240 ( .A(register__n3302), .Y(register__n11777) );
  HB1xp67_ASAP7_75t_R register___U5241 ( .A(register__n3302), .Y(register__n3301) );
  BUFx3_ASAP7_75t_R register___U5242 ( .A(register__n2854), .Y(register__n3278) );
  INVxp67_ASAP7_75t_R register___U5243 ( .A(register__n5314), .Y(register__n6724) );
  AO22x1_ASAP7_75t_R register___U5244 ( .A1(register__n9384), .A2(register__net91683), .B1(register__n9380), .B2(register__n1349), 
        .Y(register__n10874) );
  AOI22xp33_ASAP7_75t_R register___U5245 ( .A1(register__n12211), .A2(register__n1188), .B1(register__n1749), .B2(register__n1922), .Y(register__n13099) );
  CKINVDCx20_ASAP7_75t_R register___U5246 ( .A(register__n9373), .Y(register__n1749) );
  INVx2_ASAP7_75t_R register___U5247 ( .A(register__n4347), .Y(register__n7313) );
  INVxp67_ASAP7_75t_R register___U5248 ( .A(register__n2958), .Y(register__n3870) );
  HB1xp67_ASAP7_75t_R register___U5249 ( .A(register__n2959), .Y(register__n2958) );
  INVxp67_ASAP7_75t_R register___U5250 ( .A(register__n5795), .Y(register__n8672) );
  HB1xp67_ASAP7_75t_R register___U5251 ( .A(register__n12512), .Y(register__n5314) );
  INVxp67_ASAP7_75t_R register___U5252 ( .A(register__n4339), .Y(register__n6140) );
  HB1xp67_ASAP7_75t_R register___U5253 ( .A(register__n10647), .Y(register__n4339) );
  AOI22xp33_ASAP7_75t_R register___U5254 ( .A1(register__n12209), .A2(register__n587), .B1(register__n1751), .B2(register__n575), 
        .Y(register__n13222) );
  INVx1_ASAP7_75t_R register___U5255 ( .A(register__n13016), .Y(register__n1752) );
  CKINVDCx20_ASAP7_75t_R register___U5256 ( .A(register__n8767), .Y(register__n1754) );
  CKINVDCx20_ASAP7_75t_R register___U5257 ( .A(register__net90541), .Y(register__n1756) );
  HB1xp67_ASAP7_75t_R register___U5258 ( .A(register__n5443), .Y(register__n12214) );
  AOI22xp33_ASAP7_75t_R register___U5259 ( .A1(register__n10487), .A2(register__C6423_net69526), .B1(register__n10465), 
        .B2(register__net117889), .Y(register__n1757) );
  HB1xp67_ASAP7_75t_R register___U5260 ( .A(register__n13118), .Y(register__n7353) );
  AO22x1_ASAP7_75t_R register___U5261 ( .A1(register__n9802), .A2(register__n387), .B1(register__n10140), .B2(register__net120912), .Y(register__n10796) );
  AO22x1_ASAP7_75t_R register___U5262 ( .A1(register__n8757), .A2(register__net126316), .B1(register__n8083), .B2(
        net123880), .Y(register__n10625) );
  AO22x1_ASAP7_75t_R register___U5263 ( .A1(register__n8769), .A2(register__net126316), .B1(register__n10268), .B2(
        net123880), .Y(register__n10986) );
  INVx2_ASAP7_75t_R register___U5264 ( .A(register__n12213), .Y(register__n12198) );
  INVx1_ASAP7_75t_R register___U5265 ( .A(register__n11511), .Y(register__n5519) );
  HB1xp67_ASAP7_75t_R register___U5266 ( .A(register__n11380), .Y(register__n4390) );
  HB1xp67_ASAP7_75t_R register___U5267 ( .A(register__n4118), .Y(register__n4117) );
  HB1xp67_ASAP7_75t_R register___U5268 ( .A(register__n11513), .Y(register__n4118) );
  AO22x1_ASAP7_75t_R register___U5269 ( .A1(register__n9820), .A2(register__net110414), .B1(register__n10239), .B2(
        n1129), .Y(register__n11513) );
  AO22x1_ASAP7_75t_R register___U5270 ( .A1(register__n9798), .A2(register__net126316), .B1(register__n10118), .B2(
        net123880), .Y(register__n10794) );
  AO22x1_ASAP7_75t_R register___U5271 ( .A1(register__n10481), .A2(register__net126316), .B1(register__n10462), .B2(
        net123880), .Y(register__n10831) );
  AO22x1_ASAP7_75t_R register___U5272 ( .A1(register__net103558), .A2(register__net126316), .B1(register__net89553), 
        .B2(register__net123880), .Y(register__n10810) );
  AO22x1_ASAP7_75t_R register___U5273 ( .A1(register__net90689), .A2(register__n387), .B1(register__net89389), .B2(
        net120912), .Y(register__n10812) );
  AO22x1_ASAP7_75t_R register___U5274 ( .A1(register__n9720), .A2(register__net126316), .B1(register__n10160), .B2(
        net123880), .Y(register__n10647) );
  AO22x1_ASAP7_75t_R register___U5275 ( .A1(register__net114505), .A2(register__C6422_net60445), .B1(
        net112594), .B2(register__C6422_net60443), .Y(register__n11093) );
  AO22x1_ASAP7_75t_R register___U5276 ( .A1(register__n9792), .A2(register__net120789), .B1(register__n10195), .B2(
        C6422_net60443), .Y(register__n11117) );
  AO22x1_ASAP7_75t_R register___U5277 ( .A1(register__n8779), .A2(register__n38), .B1(register__n9371), .B2(
        C6422_net60443), .Y(register__n11144) );
  AO22x1_ASAP7_75t_R register___U5278 ( .A1(register__n9750), .A2(register__n38), .B1(register__n10126), .B2(
        C6422_net60443), .Y(register__n10775) );
  AO22x1_ASAP7_75t_R register___U5279 ( .A1(register__net96767), .A2(register__n38), .B1(register__net95073), .B2(
        C6422_net60443), .Y(register__n10814) );
  AO22x1_ASAP7_75t_R register___U5280 ( .A1(register__n10487), .A2(register__n38), .B1(register__n10465), .B2(
        C6422_net60443), .Y(register__n10835) );
  AO22x1_ASAP7_75t_R register___U5281 ( .A1(register__n9794), .A2(register__n38), .B1(register__n10197), .B2(
        C6422_net70678), .Y(register__n10798) );
  AO22x1_ASAP7_75t_R register___U5282 ( .A1(register__n10485), .A2(register__net126316), .B1(register__n10458), .B2(
        net123879), .Y(register__n10561) );
  AO22x1_ASAP7_75t_R register___U5283 ( .A1(register__n9268), .A2(register__C6422_net60408), .B1(register__n10191), 
        .B2(register__n834), .Y(register__n11109) );
  HB1xp67_ASAP7_75t_R register___U5284 ( .A(register__n11778), .Y(register__n11768) );
  AO22x1_ASAP7_75t_R register___U5285 ( .A1(register__n9621), .A2(register__n38), .B1(register__n10076), .B2(
        C6422_net60443), .Y(register__n10969) );
  BUFx2_ASAP7_75t_R register___U5286 ( .A(register__n5109), .Y(register__n5108) );
  AO22x1_ASAP7_75t_R register___U5287 ( .A1(register__n9736), .A2(register__net117657), .B1(register__n9319), .B2(register__n839), 
        .Y(register__n10744) );
  AOI21xp33_ASAP7_75t_R register___U5288 ( .A1(register__net110413), .A2(register__net96767), .B(register__n2716), .Y(
        n2736) );
  HB1xp67_ASAP7_75t_R register___U5289 ( .A(register__n10689), .Y(register__n5800) );
  AO22x1_ASAP7_75t_R register___U5290 ( .A1(register__n9820), .A2(register__net120789), .B1(register__n10239), .B2(
        C6422_net70678), .Y(register__n10902) );
  AO22x1_ASAP7_75t_R register___U5291 ( .A1(register__n9413), .A2(register__n1867), .B1(register__n10181), .B2(register__n91), 
        .Y(register__n10646) );
  AO22x1_ASAP7_75t_R register___U5292 ( .A1(register__n9883), .A2(register__C6422_net60415), .B1(register__n10317), 
        .B2(register__net88727), .Y(register__n10854) );
  AO22x1_ASAP7_75t_R register___U5293 ( .A1(register__n9778), .A2(register__C6422_net60445), .B1(register__n10164), 
        .B2(register__C6422_net60443), .Y(register__n10651) );
  HB1xp67_ASAP7_75t_R register___U5294 ( .A(register__n4332), .Y(register__n4331) );
  HB1xp67_ASAP7_75t_R register___U5295 ( .A(register__n10628), .Y(register__n4332) );
  AO22x1_ASAP7_75t_R register___U5296 ( .A1(register__n9260), .A2(register__C6422_net60415), .B1(register__n9923), .B2(
        net88727), .Y(register__n10628) );
  BUFx2_ASAP7_75t_R register___U5297 ( .A(register__n4111), .Y(register__n4110) );
  HB1xp67_ASAP7_75t_R register___U5298 ( .A(register__n10924), .Y(register__n4111) );
  AO22x1_ASAP7_75t_R register___U5299 ( .A1(register__n9756), .A2(register__C6422_net60415), .B1(register__n9063), .B2(
        net88727), .Y(register__n11116) );
  HB1xp67_ASAP7_75t_R register___U5300 ( .A(register__n10651), .Y(register__n5109) );
  HB1xp67_ASAP7_75t_R register___U5301 ( .A(register__n5929), .Y(register__n11833) );
  BUFx6f_ASAP7_75t_R register___U5302 ( .A(register__n3707), .Y(register__n3539) );
  BUFx6f_ASAP7_75t_R register___U5303 ( .A(register__n3539), .Y(register__n4817) );
  BUFx6f_ASAP7_75t_R register___U5304 ( .A(register__n5524), .Y(register__n11834) );
  BUFx6f_ASAP7_75t_R register___U5305 ( .A(register__n4817), .Y(register__n11912) );
  BUFx3_ASAP7_75t_R register___U5306 ( .A(register__n4818), .Y(register__n3540) );
  BUFx3_ASAP7_75t_R register___U5307 ( .A(register__n11835), .Y(register__n5044) );
  BUFx3_ASAP7_75t_R register___U5308 ( .A(register__n11835), .Y(register__n11830) );
  BUFx12f_ASAP7_75t_R register___U5309 ( .A(register__n7327), .Y(register__n11915) );
  INVx2_ASAP7_75t_R register___U5310 ( .A(register__n5471), .Y(register__n9225) );
  INVx2_ASAP7_75t_R register___U5311 ( .A(register__n5151), .Y(register__n7969) );
  BUFx3_ASAP7_75t_R register___U5312 ( .A(register__n11620), .Y(register__n5825) );
  BUFx3_ASAP7_75t_R register___U5313 ( .A(register__n7304), .Y(register__n4812) );
  INVx1_ASAP7_75t_R register___U5314 ( .A(register__n11717), .Y(register__n1761) );
  BUFx3_ASAP7_75t_R register___U5315 ( .A(register__n11302), .Y(register__n5152) );
  AO22x1_ASAP7_75t_R register___U5316 ( .A1(register__n9339), .A2(register__C6422_net60415), .B1(register__n9325), .B2(
        net88727), .Y(register__n10564) );
  NAND3xp33_ASAP7_75t_R register___U5317 ( .A(register__n11714), .B(register__n1085), .C(register__n11721), .Y(register__n1762)
         );
  CKINVDCx20_ASAP7_75t_R register___U5318 ( .A(register__net112297), .Y(register__n1763) );
  AO22x1_ASAP7_75t_R register___U5319 ( .A1(register__n8811), .A2(register__net91683), .B1(register__n8819), .B2(register__n1346), 
        .Y(register__n11046) );
  INVxp67_ASAP7_75t_R register___U5320 ( .A(register__n3966), .Y(register__n8668) );
  INVxp67_ASAP7_75t_R register___U5321 ( .A(register__n13164), .Y(register__n5938) );
  NAND2xp33_ASAP7_75t_R register___U5322 ( .A(register__n9732), .B(register__net102299), .Y(register__n1764) );
  NAND2xp33_ASAP7_75t_R register___U5323 ( .A(register__n10303), .B(register__n422), .Y(register__n1765) );
  NAND2xp33_ASAP7_75t_R register___U5324 ( .A(register__n1764), .B(register__n1765), .Y(register__n11632) );
  AND3x2_ASAP7_75t_R register___U5325 ( .A(register__n5535), .B(register__n4263), .C(register__n5536), .Y(register__n1766) );
  AND2x2_ASAP7_75t_R register___U5326 ( .A(register__n5843), .B(register__n1766), .Y(register__n11617) );
  BUFx2_ASAP7_75t_R register___U5327 ( .A(register__n5537), .Y(register__n4263) );
  BUFx12f_ASAP7_75t_R register___U5328 ( .A(register__n3938), .Y(register__n11920) );
  BUFx12f_ASAP7_75t_R register___U5329 ( .A(register__n11920), .Y(register__n11918) );
  INVx2_ASAP7_75t_R register___U5330 ( .A(register__n3422), .Y(register__n4034) );
  BUFx6f_ASAP7_75t_R register___U5331 ( .A(register__n11843), .Y(register__n4604) );
  INVx6_ASAP7_75t_R register___U5332 ( .A(register__n3735), .Y(register__n3736) );
  BUFx3_ASAP7_75t_R register___U5333 ( .A(register__n11841), .Y(register__n11919) );
  BUFx3_ASAP7_75t_R register___U5334 ( .A(register__n4603), .Y(register__n3212) );
  BUFx3_ASAP7_75t_R register___U5335 ( .A(register__n4603), .Y(register__n3384) );
  BUFx3_ASAP7_75t_R register___U5336 ( .A(register__n11841), .Y(register__n11837) );
  BUFx3_ASAP7_75t_R register___U5337 ( .A(register__n3736), .Y(register__n3216) );
  BUFx6f_ASAP7_75t_R register___U5338 ( .A(register__n4844), .Y(register__n3329) );
  BUFx6f_ASAP7_75t_R register___U5339 ( .A(register__n4844), .Y(register__n11916) );
  BUFx2_ASAP7_75t_R register___U5340 ( .A(register__n3991), .Y(register__n3422) );
  INVxp67_ASAP7_75t_R register___U5341 ( .A(register__n4202), .Y(register__n7028) );
  INVxp67_ASAP7_75t_R register___U5342 ( .A(register__n4286), .Y(register__n5843) );
  HB1xp67_ASAP7_75t_R register___U5343 ( .A(register__n4287), .Y(register__n4286) );
  BUFx6f_ASAP7_75t_R register___U5344 ( .A(register__n11818), .Y(register__n5103) );
  BUFx12f_ASAP7_75t_R register___U5345 ( .A(register__n5103), .Y(register__n3734) );
  BUFx6f_ASAP7_75t_R register___U5346 ( .A(register__n11899), .Y(register__n11897) );
  INVx1_ASAP7_75t_R register___U5347 ( .A(register__n10643), .Y(register__n7936) );
  INVxp33_ASAP7_75t_R register___U5348 ( .A(register__n10650), .Y(register__n1768) );
  HB1xp67_ASAP7_75t_R register___U5349 ( .A(register__n11632), .Y(register__n4287) );
  INVxp67_ASAP7_75t_R register___U5350 ( .A(register__n5288), .Y(register__n7639) );
  HB1xp67_ASAP7_75t_R register___U5351 ( .A(register__n5289), .Y(register__n5288) );
  AO22x1_ASAP7_75t_R register___U5352 ( .A1(register__n9881), .A2(register__C6422_net60445), .B1(register__n10321), 
        .B2(register__C6422_net60443), .Y(register__n10855) );
  INVxp67_ASAP7_75t_R register___U5353 ( .A(register__n5999), .Y(register__n7964) );
  HB1xp67_ASAP7_75t_R register___U5354 ( .A(register__n6000), .Y(register__n5999) );
  INVx1_ASAP7_75t_R register___U5355 ( .A(register__n11363), .Y(register__n1769) );
  AND2x2_ASAP7_75t_R register___U5356 ( .A(register__n8289), .B(register__n11342), .Y(register__n1770) );
  INVx1_ASAP7_75t_R register___U5357 ( .A(register__n11344), .Y(register__n8289) );
  HB1xp67_ASAP7_75t_R register___U5358 ( .A(register__n3883), .Y(register__n3882) );
  HB1xp67_ASAP7_75t_R register___U5359 ( .A(register__n12548), .Y(register__n3883) );
  HB1xp67_ASAP7_75t_R register___U5360 ( .A(register__n1768), .Y(register__n4338) );
  AO22x1_ASAP7_75t_R register___U5361 ( .A1(register__n9615), .A2(register__net126316), .B1(register__n10084), .B2(
        net123880), .Y(register__n10605) );
  AOI21xp33_ASAP7_75t_R register___U5362 ( .A1(register__C6423_net74857), .A2(register__net89565), .B(register__n2551), 
        .Y(register__n2572) );
  AO22x1_ASAP7_75t_R register___U5363 ( .A1(register__net90249), .A2(register__net93569), .B1(register__net89049), .B2(
        C6423_net74855), .Y(register__n11615) );
  HB1xp67_ASAP7_75t_R register___U5364 ( .A(register__n3967), .Y(register__n3966) );
  HB1xp67_ASAP7_75t_R register___U5365 ( .A(register__n12499), .Y(register__n1773) );
  BUFx12f_ASAP7_75t_R register___U5366 ( .A(register__n3021), .Y(register__n6720) );
  BUFx12f_ASAP7_75t_R register___U5367 ( .A(register__n6720), .Y(register__n11887) );
  HB1xp67_ASAP7_75t_R register___U5368 ( .A(register__n5504), .Y(register__n11800) );
  BUFx6f_ASAP7_75t_R register___U5369 ( .A(register__n3674), .Y(register__n2960) );
  HB1xp67_ASAP7_75t_R register___U5370 ( .A(register__n5501), .Y(register__n11802) );
  INVxp33_ASAP7_75t_R register___U5371 ( .A(register__n1646), .Y(register__n1775) );
  INVx1_ASAP7_75t_R register___U5372 ( .A(register__n1785), .Y(register__n1786) );
  HB1xp67_ASAP7_75t_R register___U5373 ( .A(register__n10855), .Y(register__n5289) );
  AO22x1_ASAP7_75t_R register___U5374 ( .A1(register__n8775), .A2(register__n38), .B1(register__n10144), .B2(
        C6422_net60443), .Y(register__n10751) );
  AO22x1_ASAP7_75t_R register___U5375 ( .A1(register__n9623), .A2(register__n38), .B1(register__n7487), .B2(
        C6422_net60443), .Y(register__n10925) );
  AO22x1_ASAP7_75t_R register___U5376 ( .A1(register__net93508), .A2(register__C6422_net60445), .B1(register__net93420), 
        .B2(register__C6422_net60443), .Y(register__n11009) );
  AO22x1_ASAP7_75t_R register___U5377 ( .A1(register__n9830), .A2(register__n38), .B1(register__n10271), .B2(
        C6422_net60443), .Y(register__n10990) );
  BUFx6f_ASAP7_75t_R register___U5378 ( .A(register__n3674), .Y(register__n3546) );
  INVx1_ASAP7_75t_R register___U5379 ( .A(register__n10773), .Y(register__n6829) );
  HB1xp67_ASAP7_75t_R register___U5380 ( .A(register__n12527), .Y(register__n5973) );
  HB1xp67_ASAP7_75t_R register___U5381 ( .A(register__n12523), .Y(register__n4526) );
  AO22x1_ASAP7_75t_R register___U5382 ( .A1(register__n9668), .A2(register__C6422_net60415), .B1(register__n9915), .B2(
        net88727), .Y(register__n10968) );
  BUFx3_ASAP7_75t_R register___U5383 ( .A(register__n10834), .Y(register__n4022) );
  AO22x1_ASAP7_75t_R register___U5384 ( .A1(register__n9303), .A2(register__C6422_net60415), .B1(register__n6949), .B2(
        net88727), .Y(register__n10901) );
  AO22x1_ASAP7_75t_R register___U5385 ( .A1(register__n9672), .A2(register__C6422_net60415), .B1(register__n9919), .B2(
        net88727), .Y(register__n10924) );
  HB1xp67_ASAP7_75t_R register___U5386 ( .A(register__n12843), .Y(register__n4666) );
  HB1xp67_ASAP7_75t_R register___U5387 ( .A(register__n12844), .Y(register__n7123) );
  HB1xp67_ASAP7_75t_R register___U5388 ( .A(register__n11243), .Y(register__n6000) );
  AO22x1_ASAP7_75t_R register___U5389 ( .A1(register__n9780), .A2(register__n387), .B1(register__n10096), .B2(register__net120912), .Y(register__n10649) );
  OAI22xp5_ASAP7_75t_R register___U5390 ( .A1(register__n54), .A2(register__n7939), .B1(register__net61369), .B2(register__n12094), .Y(read_reg_data_1[9]) );
  AOI22xp33_ASAP7_75t_R register___U5391 ( .A1(register__net63376), .A2(register__n1622), .B1(register__n1799), .B2(
        n1647), .Y(register__n12754) );
  CKINVDCx20_ASAP7_75t_R register___U5392 ( .A(register__n10263), .Y(register__n1799) );
  INVxp67_ASAP7_75t_R register___U5393 ( .A(register__n3010), .Y(register__n6195) );
  AO22x1_ASAP7_75t_R register___U5394 ( .A1(register__net88472), .A2(register__net121619), .B1(register__net119537), 
        .B2(register__net126625), .Y(register__n11011) );
  INVx1_ASAP7_75t_R register___U5395 ( .A(register__n10749), .Y(register__n1804) );
  AND2x2_ASAP7_75t_R register___U5396 ( .A(register__n10734), .B(register__n10732), .Y(register__n1805) );
  AND3x1_ASAP7_75t_R register___U5397 ( .A(register__n1805), .B(register__n10733), .C(register__n771), .Y(register__n9179) );
  AND2x2_ASAP7_75t_R register___U5398 ( .A(register__n1806), .B(register__n1882), .Y(register__n10679) );
  HB1xp67_ASAP7_75t_R register___U5399 ( .A(register__n12551), .Y(register__n4201) );
  INVxp33_ASAP7_75t_R register___U5400 ( .A(register__n7633), .Y(register__n1812) );
  INVxp33_ASAP7_75t_R register___U5401 ( .A(register__n5516), .Y(register__n1823) );
  INVxp67_ASAP7_75t_R register___U5402 ( .A(register__n1825), .Y(register__n1826) );
  INVxp67_ASAP7_75t_R register___U5403 ( .A(register__n1829), .Y(register__n1830) );
  INVx2_ASAP7_75t_R register___U5404 ( .A(register__n3168), .Y(register__n1831) );
  INVx1_ASAP7_75t_R register___U5405 ( .A(register__n1831), .Y(register__n1832) );
  BUFx6f_ASAP7_75t_R register___U5406 ( .A(register__n3709), .Y(register__n9379) );
  HB1xp67_ASAP7_75t_R register___U5407 ( .A(register__n4869), .Y(register__n4868) );
  HB1xp67_ASAP7_75t_R register___U5408 ( .A(register__n12840), .Y(register__n4869) );
  HB1xp67_ASAP7_75t_R register___U5409 ( .A(register__n7119), .Y(register__n7118) );
  HB1xp67_ASAP7_75t_R register___U5410 ( .A(register__n12839), .Y(register__n7119) );
  INVxp67_ASAP7_75t_R register___U5411 ( .A(register__n5068), .Y(register__n7728) );
  HB1xp67_ASAP7_75t_R register___U5412 ( .A(register__n5069), .Y(register__n5068) );
  HB1xp67_ASAP7_75t_R register___U5413 ( .A(register__n11146), .Y(register__n5069) );
  AO22x1_ASAP7_75t_R register___U5414 ( .A1(register__n9861), .A2(register__net121619), .B1(register__n10295), .B2(
        net126625), .Y(register__n11146) );
  AO22x1_ASAP7_75t_R register___U5415 ( .A1(register__n9297), .A2(register__n930), .B1(register__n10187), .B2(register__net150894), .Y(register__n11317) );
  NOR2xp67_ASAP7_75t_R register___U5416 ( .A(register__net109880), .B(register__n1800), .Y(register__n2425) );
  INVx1_ASAP7_75t_R register___U5417 ( .A(register__n11450), .Y(register__n8751) );
  INVxp67_ASAP7_75t_R register___U5418 ( .A(register__n5799), .Y(register__n7603) );
  HB1xp67_ASAP7_75t_R register___U5419 ( .A(register__n5800), .Y(register__n5799) );
  AO22x1_ASAP7_75t_R register___U5420 ( .A1(register__n9722), .A2(register__net117658), .B1(register__n10162), .B2(register__n838), .Y(register__n10643) );
  INVxp67_ASAP7_75t_R register___U5421 ( .A(register__n4616), .Y(register__n8626) );
  HB1xp67_ASAP7_75t_R register___U5422 ( .A(register__n4617), .Y(register__n4616) );
  INVxp67_ASAP7_75t_R register___U5423 ( .A(register__n4200), .Y(register__n6169) );
  HB1xp67_ASAP7_75t_R register___U5424 ( .A(register__n4201), .Y(register__n4200) );
  BUFx12f_ASAP7_75t_R register___U5425 ( .A(register__n11918), .Y(register__n11917) );
  AO22x1_ASAP7_75t_R register___U5426 ( .A1(register__n9828), .A2(register__C6423_net74825), .B1(register__n10243), 
        .B2(register__C6423_net74851), .Y(register__n11515) );
  INVx2_ASAP7_75t_R register___U5427 ( .A(register__n11515), .Y(register__n2924) );
  AO22x1_ASAP7_75t_R register___U5428 ( .A1(register__n7555), .A2(register__n1771), .B1(register__n5877), .B2(register__net126625), .Y(register__n10695) );
  HB1xp67_ASAP7_75t_R register___U5429 ( .A(register__n5516), .Y(register__n4955) );
  AO22x1_ASAP7_75t_R register___U5430 ( .A1(register__n9274), .A2(register__C6422_net60415), .B1(register__n10263), 
        .B2(register__net88727), .Y(register__n10989) );
  AO22x1_ASAP7_75t_R register___U5431 ( .A1(register__net90401), .A2(register__C6422_net60415), .B1(register__net115976), .B2(register__net88727), .Y(register__n10711) );
  HB1xp67_ASAP7_75t_R register___U5432 ( .A(register__net109643), .Y(register__net126596) );
  BUFx12f_ASAP7_75t_R register___U5433 ( .A(register__C6422_net60401), .Y(register__net126602) );
  INVxp67_ASAP7_75t_R register___U5434 ( .A(register__n3106), .Y(register__n7321) );
  HB1xp67_ASAP7_75t_R register___U5435 ( .A(register__n3107), .Y(register__n3106) );
  AO22x1_ASAP7_75t_R register___U5436 ( .A1(register__n9710), .A2(register__net131160), .B1(register__n10040), .B2(
        net120912), .Y(register__n10833) );
  AO22x1_ASAP7_75t_R register___U5437 ( .A1(register__n7392), .A2(register__C6422_net60405), .B1(register__n4961), .B2(
        C6422_net60401), .Y(register__n11133) );
  AO22x1_ASAP7_75t_R register___U5438 ( .A1(register__n6098), .A2(register__net117658), .B1(register__n10124), .B2(register__n838), .Y(register__n10767) );
  NOR2xp67_ASAP7_75t_R register___U5439 ( .A(register__C6423_net61114), .B(register__n1691), .Y(register__n2639) );
  AO22x1_ASAP7_75t_R register___U5440 ( .A1(register__n7192), .A2(register__net126316), .B1(register__n10273), .B2(
        net123880), .Y(register__n10689) );
  HB1xp67_ASAP7_75t_R register___U5441 ( .A(register__n3011), .Y(register__n3010) );
  INVxp33_ASAP7_75t_R register___U5442 ( .A(register__n5797), .Y(register__n7601) );
  HB1xp67_ASAP7_75t_R register___U5443 ( .A(register__n10685), .Y(register__n3107) );
  INVx2_ASAP7_75t_R register___U5444 ( .A(register__n4150), .Y(register__n5385) );
  BUFx3_ASAP7_75t_R register___U5445 ( .A(register__n4151), .Y(register__n4150) );
  HB1xp67_ASAP7_75t_R register___U5446 ( .A(register__n11133), .Y(register__n2894) );
  HB1xp67_ASAP7_75t_R register___U5447 ( .A(register__n12755), .Y(register__n3608) );
  AO22x1_ASAP7_75t_R register___U5448 ( .A1(register__net117710), .A2(register__net118635), .B1(register__net89285), 
        .B2(register__net126625), .Y(register__n10714) );
  INVxp67_ASAP7_75t_R register___U5449 ( .A(register__n3886), .Y(register__n8648) );
  AO22x1_ASAP7_75t_R register___U5450 ( .A1(register__n9301), .A2(register__n929), .B1(register__n10337), .B2(register__n769), 
        .Y(register__n11675) );
  HB1xp67_ASAP7_75t_R register___U5451 ( .A(register__n9408), .Y(register__n5735) );
  AO22x1_ASAP7_75t_R register___U5452 ( .A1(register__n9696), .A2(register__C6423_net61340), .B1(register__n9967), .B2(
        n334), .Y(register__n11167) );
  AO22x1_ASAP7_75t_R register___U5453 ( .A1(register__n10497), .A2(register__C6423_net61340), .B1(register__n8787), 
        .B2(register__n334), .Y(register__n11189) );
  HB1xp67_ASAP7_75t_R register___U5454 ( .A(register__n7601), .Y(register__n5798) );
  HB1xp67_ASAP7_75t_R register___U5455 ( .A(register__n11011), .Y(register__n4617) );
  AO22x1_ASAP7_75t_R register___U5456 ( .A1(register__n5644), .A2(register__n1771), .B1(register__n6038), .B2(
        C6422_net70534), .Y(register__n10586) );
  AO22x1_ASAP7_75t_R register___U5457 ( .A1(register__net90637), .A2(register__C6423_net61340), .B1(register__net89649), 
        .B2(register__net125365), .Y(register__n11610) );
  HB1xp67_ASAP7_75t_R register___U5458 ( .A(register__n10721), .Y(register__n3011) );
  AO22x1_ASAP7_75t_R register___U5459 ( .A1(register__net93817), .A2(register__net117658), .B1(register__net89585), 
        .B2(register__n842), .Y(register__n10721) );
  HB1xp67_ASAP7_75t_R register___U5460 ( .A(register__n3887), .Y(register__n3886) );
  BUFx3_ASAP7_75t_R register___U5461 ( .A(register__n11642), .Y(register__n6029) );
  OAI22xp33_ASAP7_75t_R register___U5462 ( .A1(register__net99872), .A2(register__n2605), .B1(register__n1903), .B2(
        n2603), .Y(register__n2588) );
  INVx2_ASAP7_75t_R register___U5463 ( .A(register__n4928), .Y(register__n7956) );
  NOR2xp33_ASAP7_75t_R register___U5464 ( .A(register__n2013), .B(register__n7695), .Y(register__n1837) );
  NOR2xp33_ASAP7_75t_R register___U5465 ( .A(register__net130175), .B(register__n11664), .Y(register__n1838) );
  NOR2xp33_ASAP7_75t_R register___U5466 ( .A(register__n1837), .B(register__n1838), .Y(register__n11662) );
  BUFx2_ASAP7_75t_R register___U5467 ( .A(register__n11563), .Y(register__n5315) );
  OAI21xp33_ASAP7_75t_R register___U5468 ( .A1(register__n1800), .A2(register__n2492), .B(register__n2511), .Y(register__n2510)
         );
  HB1xp67_ASAP7_75t_R register___U5469 ( .A(register__n4706), .Y(register__n4705) );
  INVxp67_ASAP7_75t_R register___U5470 ( .A(register__n4128), .Y(register__n6176) );
  HB1xp67_ASAP7_75t_R register___U5471 ( .A(register__n4129), .Y(register__n4128) );
  NOR2xp67_ASAP7_75t_R register___U5472 ( .A(register__net103300), .B(register__n802), .Y(register__n2324) );
  INVx1_ASAP7_75t_R register___U5473 ( .A(register__n13202), .Y(register__n1839) );
  AO22x1_ASAP7_75t_R register___U5474 ( .A1(register__n9349), .A2(register__net141083), .B1(register__n9367), .B2(register__n334), 
        .Y(register__n11671) );
  NAND2xp33_ASAP7_75t_R register___U5475 ( .A(register__net90717), .B(register__C6422_net70498), .Y(register__n1840) );
  BUFx6f_ASAP7_75t_R register___U5476 ( .A(register__net89590), .Y(register__net89589) );
  INVxp67_ASAP7_75t_R register___U5477 ( .A(register__n4291), .Y(register__n5931) );
  AND3x1_ASAP7_75t_R register___U5478 ( .A(register__n267), .B(register__n63), .C(register__n7913), .Y(register__n2777) );
  HB1xp67_ASAP7_75t_R register___U5479 ( .A(register__n12773), .Y(register__n3887) );
  INVxp67_ASAP7_75t_R register___U5480 ( .A(register__n13388), .Y(read_reg_data_1[15]) );
  BUFx3_ASAP7_75t_R register___U5481 ( .A(register__n10660), .Y(register__n4929) );
  AO22x1_ASAP7_75t_R register___U5482 ( .A1(register__n9766), .A2(register__C6423_net61340), .B1(register__n10114), 
        .B2(register__net125365), .Y(register__n11631) );
  BUFx6f_ASAP7_75t_R register___U5483 ( .A(register__net107120), .Y(register__net107119) );
  AND4x1_ASAP7_75t_R register___U5484 ( .A(register__n8636), .B(register__n1556), .C(register__n5304), .D(register__n5563), .Y(
        n10779) );
  HB1xp67_ASAP7_75t_R register___U5485 ( .A(register__n12774), .Y(register__n4129) );
  HB1xp67_ASAP7_75t_R register___U5486 ( .A(register__n11510), .Y(register__n4706) );
  AO22x1_ASAP7_75t_R register___U5487 ( .A1(register__n9688), .A2(register__net123861), .B1(register__n9959), .B2(
        net125365), .Y(register__n11487) );
  HB1xp67_ASAP7_75t_R register___U5488 ( .A(register__n11189), .Y(register__n5415) );
  AO22x1_ASAP7_75t_R register___U5489 ( .A1(register__n8771), .A2(register__C6423_net61340), .B1(register__n7140), .B2(
        C6423_net69198), .Y(register__n11465) );
  AOI22xp33_ASAP7_75t_R register___U5490 ( .A1(register__n9585), .A2(register__net118635), .B1(register__n10006), .B2(
        C6422_net70534), .Y(register__n1842) );
  AO22x1_ASAP7_75t_R register___U5491 ( .A1(register__n9589), .A2(register__net121619), .B1(register__n10010), .B2(
        net126625), .Y(register__n10631) );
  AND2x2_ASAP7_75t_R register___U5492 ( .A(register__n11720), .B(register__n1953), .Y(register__n1967) );
  INVx2_ASAP7_75t_R register___U5493 ( .A(register__n11736), .Y(register__n11853) );
  INVx3_ASAP7_75t_R register___U5494 ( .A(register__n1901), .Y(register__n11735) );
  BUFx3_ASAP7_75t_R register___U5495 ( .A(register__n11735), .Y(register__n3866) );
  BUFx3_ASAP7_75t_R register___U5496 ( .A(register__n11735), .Y(register__n3867) );
  BUFx3_ASAP7_75t_R register___U5497 ( .A(register__n11735), .Y(register__n3868) );
  INVx3_ASAP7_75t_R register___U5498 ( .A(register__n2945), .Y(register__n11736) );
  AO22x1_ASAP7_75t_R register___U5499 ( .A1(register__n9351), .A2(register__n2), .B1(register__n8354), .B2(
        C6422_net60443), .Y(register__n11051) );
  INVxp67_ASAP7_75t_R register___U5500 ( .A(register__n4084), .Y(register__n5944) );
  AO22x1_ASAP7_75t_R register___U5501 ( .A1(register__n9726), .A2(register__net109204), .B1(register__n5680), .B2(register__n59), 
        .Y(register__n10650) );
  AO22x1_ASAP7_75t_R register___U5502 ( .A1(register__n9901), .A2(register__n1771), .B1(register__n10333), .B2(
        net126625), .Y(register__n11076) );
  AO22x1_ASAP7_75t_R register___U5503 ( .A1(register__n8777), .A2(register__C6423_net61340), .B1(register__n10112), 
        .B2(register__net125365), .Y(register__n11510) );
  INVxp67_ASAP7_75t_R register___U5504 ( .A(register__n4523), .Y(register__n6129) );
  AO22x1_ASAP7_75t_R register___U5505 ( .A1(register__n9738), .A2(register__n387), .B1(register__n10305), .B2(register__net120912), .Y(register__n10749) );
  AO22x1_ASAP7_75t_R register___U5506 ( .A1(register__n9341), .A2(register__net117658), .B1(register__n8351), .B2(register__n837), 
        .Y(register__n10685) );
  AND3x1_ASAP7_75t_R register___U5507 ( .A(register__n7914), .B(register__n7915), .C(register__n7600), .Y(register__n2788) );
  AO22x1_ASAP7_75t_R register___U5508 ( .A1(register__n9611), .A2(register__C6423_net61343), .B1(register__n10078), 
        .B2(register__net129787), .Y(register__n11532) );
  AO22x1_ASAP7_75t_R register___U5509 ( .A1(register__n9770), .A2(register__C6423_net61343), .B1(register__n10120), 
        .B2(register__net129787), .Y(register__n11464) );
  AO22x1_ASAP7_75t_R register___U5510 ( .A1(register__n6838), .A2(register__C6423_net61343), .B1(register__n10072), 
        .B2(register__net122313), .Y(register__n11572) );
  AO22x1_ASAP7_75t_R register___U5511 ( .A1(register__n9720), .A2(register__C6423_net61343), .B1(register__n10160), 
        .B2(register__net129787), .Y(register__n11312) );
  AO22x1_ASAP7_75t_R register___U5512 ( .A1(register__n9609), .A2(register__C6423_net61343), .B1(register__n10074), 
        .B2(register__C6423_net69272), .Y(register__n11553) );
  HB1xp67_ASAP7_75t_R register___U5513 ( .A(register__n12514), .Y(register__n6760) );
  HB1xp67_ASAP7_75t_R register___U5514 ( .A(register__n10692), .Y(register__n5797) );
  BUFx3_ASAP7_75t_R register___U5515 ( .A(register__n11420), .Y(register__n5424) );
  BUFx12f_ASAP7_75t_R register___U5516 ( .A(register__net126602), .Y(register__net126601) );
  INVxp67_ASAP7_75t_R register___U5517 ( .A(register__n2876), .Y(register__n3996) );
  INVxp67_ASAP7_75t_R register___U5518 ( .A(register__n4246), .Y(register__n5522) );
  HB1xp67_ASAP7_75t_R register___U5519 ( .A(register__n10726), .Y(register__n4246) );
  HB1xp67_ASAP7_75t_R register___U5520 ( .A(register__n11140), .Y(register__n4819) );
  OAI22xp33_ASAP7_75t_R register___U5521 ( .A1(register__n6679), .A2(register__n954), .B1(register__n10440), .B2(register__n959), 
        .Y(register__n1855) );
  CKINVDCx20_ASAP7_75t_R register___U5522 ( .A(register__net95244), .Y(register__n1856) );
  CKINVDCx20_ASAP7_75t_R register___U5523 ( .A(register__net98849), .Y(register__n1857) );
  INVxp67_ASAP7_75t_R register___U5524 ( .A(register__n4304), .Y(register__n6685) );
  AND3x1_ASAP7_75t_R register___U5525 ( .A(register__n9396), .B(register__n1842), .C(register__n8266), .Y(register__n2779) );
  HB1xp67_ASAP7_75t_R register___U5526 ( .A(register__n2877), .Y(register__n2876) );
  AO22x1_ASAP7_75t_R register___U5527 ( .A1(register__n8777), .A2(register__net129747), .B1(register__n10112), .B2(
        net123857), .Y(register__n10899) );
  AO22x1_ASAP7_75t_R register___U5528 ( .A1(register__n8771), .A2(register__n1853), .B1(register__n7141), .B2(register__net139537), .Y(register__n10852) );
  HB1xp67_ASAP7_75t_R register___U5529 ( .A(register__n4524), .Y(register__n4523) );
  HB1xp67_ASAP7_75t_R register___U5530 ( .A(register__n13313), .Y(register__n4524) );
  HB1xp67_ASAP7_75t_R register___U5531 ( .A(register__n4085), .Y(register__n4084) );
  AO22x1_ASAP7_75t_R register___U5532 ( .A1(register__n9290), .A2(register__net122579), .B1(register__n9937), .B2(
        net150889), .Y(register__n11257) );
  AO22x1_ASAP7_75t_R register___U5533 ( .A1(register__n6957), .A2(register__net122579), .B1(register__n10471), .B2(
        net150896), .Y(register__n11514) );
  INVx1_ASAP7_75t_R register___U5534 ( .A(register__n10895), .Y(register__n1858) );
  CKINVDCx20_ASAP7_75t_R register___U5535 ( .A(register__n9421), .Y(register__n1860) );
  HB1xp67_ASAP7_75t_R register___U5536 ( .A(register__n4305), .Y(register__n4304) );
  INVxp67_ASAP7_75t_R register___U5537 ( .A(register__n6495), .Y(register__n8037) );
  HB1xp67_ASAP7_75t_R register___U5538 ( .A(register__n6496), .Y(register__n6495) );
  AOI22xp33_ASAP7_75t_R register___U5539 ( .A1(register__net64054), .A2(register__n470), .B1(register__n1862), .B2(register__n460), .Y(register__n12934) );
  CKINVDCx20_ASAP7_75t_R register___U5540 ( .A(register__net89401), .Y(register__n1862) );
  INVx2_ASAP7_75t_R register___U5541 ( .A(register__net64042), .Y(register__net64008) );
  BUFx3_ASAP7_75t_R register___U5542 ( .A(register__net104773), .Y(register__n1863) );
  INVx2_ASAP7_75t_R register___U5543 ( .A(register__net104772), .Y(register__n1865) );
  BUFx6f_ASAP7_75t_R register___U5544 ( .A(register__net91683), .Y(register__net104773) );
  BUFx6f_ASAP7_75t_R register___U5545 ( .A(register__net137523), .Y(register__net137521) );
  CKINVDCx20_ASAP7_75t_R register___U5546 ( .A(register__n8761), .Y(register__n1868) );
  CKINVDCx20_ASAP7_75t_R register___U5547 ( .A(register__n9947), .Y(register__n1869) );
  INVx1_ASAP7_75t_R register___U5548 ( .A(register__n13043), .Y(register__n1870) );
  OAI22xp33_ASAP7_75t_R register___U5549 ( .A1(register__net62828), .A2(register__n892), .B1(register__net90233), .B2(
        n902), .Y(register__n1871) );
  AO22x1_ASAP7_75t_R register___U5550 ( .A1(register__n9599), .A2(register__n39), .B1(register__n10022), .B2(
        C6422_net60399), .Y(register__n10829) );
  AO22x1_ASAP7_75t_R register___U5551 ( .A1(register__net95344), .A2(register__n39), .B1(register__net88512), .B2(
        C6422_net60399), .Y(register__n10723) );
  INVxp67_ASAP7_75t_R register___U5552 ( .A(register__n3828), .Y(register__n5218) );
  AND3x2_ASAP7_75t_R register___U5553 ( .A(register__n731), .B(register__n11714), .C(rs2[0]), .Y(
        n11719) );
  AO22x1_ASAP7_75t_R register___U5554 ( .A1(register__net90673), .A2(register__n1853), .B1(register__net89661), .B2(
        net123857), .Y(register__n10726) );
  AO22x1_ASAP7_75t_R register___U5555 ( .A1(register__n7574), .A2(register__net109204), .B1(register__n10297), .B2(register__n59), 
        .Y(register__n11140) );
  INVxp33_ASAP7_75t_R register___U5556 ( .A(register__net137463), .Y(register__n1873) );
  INVxp67_ASAP7_75t_R register___U5557 ( .A(register__n5093), .Y(register__n6692) );
  HB1xp67_ASAP7_75t_R register___U5558 ( .A(register__n5094), .Y(register__n5093) );
  HB1xp67_ASAP7_75t_R register___U5559 ( .A(register__n10705), .Y(register__n2877) );
  AO22x1_ASAP7_75t_R register___U5560 ( .A1(register__net90393), .A2(register__n413), .B1(register__net89277), .B2(
        net126602), .Y(register__n10705) );
  HB1xp67_ASAP7_75t_R register___U5561 ( .A(register__n10727), .Y(register__n6496) );
  HB1xp67_ASAP7_75t_R register___U5562 ( .A(register__n13250), .Y(register__n4305) );
  AO22x1_ASAP7_75t_R register___U5563 ( .A1(register__n9722), .A2(register__net128121), .B1(register__n10162), .B2(
        n1999), .Y(register__n11308) );
  INVxp67_ASAP7_75t_R register___U5564 ( .A(register__n3142), .Y(register__n7599) );
  HB1xp67_ASAP7_75t_R register___U5565 ( .A(register__n3143), .Y(register__n3142) );
  HB1xp67_ASAP7_75t_R register___U5566 ( .A(register__n13055), .Y(register__n5094) );
  INVx1_ASAP7_75t_R register___U5567 ( .A(register__n11611), .Y(register__n1874) );
  AO22x1_ASAP7_75t_R register___U5568 ( .A1(register__n9879), .A2(register__n482), .B1(register__n10157), .B2(
        C6423_net61348), .Y(register__n11385) );
  AO22x1_ASAP7_75t_R register___U5569 ( .A1(register__n9652), .A2(register__net109849), .B1(register__n9979), .B2(register__n649), 
        .Y(register__n11239) );
  AO22x1_ASAP7_75t_R register___U5570 ( .A1(register__n481), .A2(register__n9744), .B1(register__n10132), .B2(register__n644), 
        .Y(register__n11405) );
  NOR2xp67_ASAP7_75t_R register___U5571 ( .A(register__n_cell_124938_net165675), .B(register__n2469), .Y(
        n2471) );
  HB1xp67_ASAP7_75t_R register___U5572 ( .A(register__n3829), .Y(register__n3828) );
  HB1xp67_ASAP7_75t_R register___U5573 ( .A(register__n13038), .Y(register__n3829) );
  INVx1_ASAP7_75t_R register___U5574 ( .A(register__n13267), .Y(register__n1875) );
  HB1xp67_ASAP7_75t_R register___U5575 ( .A(register__n11609), .Y(register__n7064) );
  CKINVDCx20_ASAP7_75t_R register___U5576 ( .A(register__net93508), .Y(register__n1877) );
  HB1xp67_ASAP7_75t_R register___U5577 ( .A(register__n2833), .Y(register__n2832) );
  HB1xp67_ASAP7_75t_R register___U5578 ( .A(register__n10828), .Y(register__n2833) );
  INVxp67_ASAP7_75t_R register___U5579 ( .A(register__n2832), .Y(register__n3699) );
  HB1xp67_ASAP7_75t_R register___U5580 ( .A(register__n7945), .Y(register__n3634) );
  INVxp33_ASAP7_75t_R register___U5581 ( .A(register__n3632), .Y(register__n7945) );
  AO22x1_ASAP7_75t_R register___U5582 ( .A1(register__n7823), .A2(register__net146144), .B1(register__n8506), .B2(
        net126601), .Y(register__n10895) );
  AO22x2_ASAP7_75t_R register___U5583 ( .A1(register__net63216), .A2(register__n673), .B1(register__C6423_net61141), 
        .B2(register__n701), .Y(register__n1878) );
  INVx1_ASAP7_75t_R register___U5584 ( .A(register__n12806), .Y(register__n1879) );
  AO22x1_ASAP7_75t_R register___U5585 ( .A1(register__n9712), .A2(register__n85), .B1(register__n10042), .B2(
        C6423_net61335), .Y(register__n11335) );
  HB1xp67_ASAP7_75t_R register___U5586 ( .A(register__n2157), .Y(register__C6423_net60474) );
  HB1xp67_ASAP7_75t_R register___U5587 ( .A(register__n6198), .Y(register__n3130) );
  INVxp33_ASAP7_75t_R register___U5588 ( .A(register__n3129), .Y(register__n6198) );
  AND2x2_ASAP7_75t_R register___U5589 ( .A(register__n1040), .B(register__n10678), .Y(register__n1881) );
  INVxp67_ASAP7_75t_R register___U5590 ( .A(register__n5008), .Y(register__n7079) );
  HB1xp67_ASAP7_75t_R register___U5591 ( .A(register__n13312), .Y(register__n5008) );
  INVxp67_ASAP7_75t_R register___U5592 ( .A(register__n12805), .Y(register__n6744) );
  HB1xp67_ASAP7_75t_R register___U5593 ( .A(register__n3342), .Y(register__n12382) );
  AO22x1_ASAP7_75t_R register___U5594 ( .A1(register__n8930), .A2(register__n85), .B1(register__n10038), .B2(register__n422), .Y(
        n11488) );
  AO22x1_ASAP7_75t_R register___U5595 ( .A1(register__n9738), .A2(register__net129017), .B1(register__n10305), .B2(
        C6423_net61335), .Y(register__n11380) );
  AO22x1_ASAP7_75t_R register___U5596 ( .A1(register__n9857), .A2(register__net102299), .B1(register__n10327), .B2(register__n422), .Y(register__n11717) );
  BUFx12f_ASAP7_75t_R register___U5597 ( .A(register__n1880), .Y(register__n12386) );
  INVx6_ASAP7_75t_R register___U5598 ( .A(register__n12386), .Y(register__n12371) );
  AOI21xp33_ASAP7_75t_R register___U5599 ( .A1(register__C6423_net68948), .A2(register__net93639), .B(register__n1902), 
        .Y(register__n2721) );
  AO22x1_ASAP7_75t_R register___U5600 ( .A1(register__n10477), .A2(register__C6423_net61326), .B1(register__n10456), 
        .B2(register__n2137), .Y(register__n11329) );
  AO22x1_ASAP7_75t_R register___U5601 ( .A1(register__n9734), .A2(register__net128122), .B1(register__n8510), .B2(register__n2000), .Y(register__n11588) );
  AO22x1_ASAP7_75t_R register___U5602 ( .A1(register__n9270), .A2(register__net128122), .B1(register__n10193), .B2(
        n2001), .Y(register__n11416) );
  AO22x1_ASAP7_75t_R register___U5603 ( .A1(register__n9341), .A2(register__net124706), .B1(register__n8351), .B2(register__n2001), .Y(register__n11354) );
  AO22x1_ASAP7_75t_R register___U5604 ( .A1(register__net93793), .A2(register__C6423_net61326), .B1(register__net103569), .B2(register__net120961), .Y(register__n11606) );
  INVxp67_ASAP7_75t_R register___U5605 ( .A(register__n3964), .Y(register__n6167) );
  HB1xp67_ASAP7_75t_R register___U5606 ( .A(register__n3965), .Y(register__n3964) );
  AO22x1_ASAP7_75t_R register___U5607 ( .A1(register__net90541), .A2(register__net137440), .B1(register__net112345), 
        .B2(register__net125803), .Y(register__n11609) );
  HB1xp67_ASAP7_75t_R register___U5608 ( .A(register__n13247), .Y(register__n4209) );
  NOR2xp67_ASAP7_75t_R register___U5609 ( .A(register__n1800), .B(register__n2530), .Y(register__n2534) );
  NOR2xp67_ASAP7_75t_R register___U5610 ( .A(register__net107836), .B(register__n1800), .Y(register__n2591) );
  AO22x1_ASAP7_75t_R register___U5611 ( .A1(register__net90257), .A2(register__n85), .B1(register__net89645), .B2(register__n422), 
        .Y(register__n11611) );
  HB1xp67_ASAP7_75t_R register___U5612 ( .A(register__n3633), .Y(register__n3632) );
  HB1xp67_ASAP7_75t_R register___U5613 ( .A(register__n10792), .Y(register__n3633) );
  HB1xp67_ASAP7_75t_R register___U5614 ( .A(register__n12927), .Y(register__n3685) );
  BUFx5_ASAP7_75t_R register___U5615 ( .A(register__n1153), .Y(register__n12381) );
  BUFx3_ASAP7_75t_R register___U5616 ( .A(register__n780), .Y(register__n3199) );
  INVxp67_ASAP7_75t_R register___U5617 ( .A(register__n3970), .Y(register__n6136) );
  HB1xp67_ASAP7_75t_R register___U5618 ( .A(register__n12939), .Y(register__n3970) );
  CKINVDCx20_ASAP7_75t_R register___U5619 ( .A(register__n9638), .Y(register__n1883) );
  HB1xp67_ASAP7_75t_R register___U5620 ( .A(register__n4292), .Y(register__n4291) );
  INVxp67_ASAP7_75t_R register___U5621 ( .A(register__n13083), .Y(register__n7950) );
  AO22x1_ASAP7_75t_R register___U5622 ( .A1(register__n9842), .A2(register__net121619), .B1(register__n10267), .B2(
        net126625), .Y(register__n11053) );
  AO22x1_ASAP7_75t_R register___U5623 ( .A1(register__net90529), .A2(register__net118635), .B1(register__net89405), 
        .B2(register__net126625), .Y(register__n10816) );
  INVxp33_ASAP7_75t_R register___U5624 ( .A(register__n12214), .Y(register__n3759) );
  INVxp67_ASAP7_75t_R register___U5625 ( .A(register__n3174), .Y(register__n5543) );
  HB1xp67_ASAP7_75t_R register___U5626 ( .A(register__n12908), .Y(register__n3174) );
  AOI21xp33_ASAP7_75t_R register___U5627 ( .A1(register__n1074), .A2(register__net89581), .B(register__n2612), .Y(register__n2632) );
  AO22x1_ASAP7_75t_R register___U5628 ( .A1(register__n9792), .A2(register__net110414), .B1(register__n10195), .B2(
        n1129), .Y(register__n11696) );
  NAND2xp67_ASAP7_75t_R register___U5629 ( .A(register__net128109), .B(register__net90925), .Y(register__n2453) );
  NOR3x1_ASAP7_75t_R register___U5630 ( .A(register__n10782), .B(register__n2254), .C(register__n2253), .Y(register__n7273) );
  HB1xp67_ASAP7_75t_R register___U5631 ( .A(register__n12546), .Y(register__n4292) );
  HB1xp67_ASAP7_75t_R register___U5632 ( .A(register__n1282), .Y(register__n1884) );
  HB1xp67_ASAP7_75t_R register___U5633 ( .A(register__n2310), .Y(register__n1885) );
  BUFx4f_ASAP7_75t_R register___U5634 ( .A(register__n2584), .Y(register__n2559) );
  INVx4_ASAP7_75t_R register___U5635 ( .A(register__n2559), .Y(register__n1886) );
  OR2x2_ASAP7_75t_R register___U5636 ( .A(register__net109215), .B(register__n1684), .Y(register__n2312) );
  INVx2_ASAP7_75t_R register___U5637 ( .A(register__n2312), .Y(register__n1888) );
  NOR2x1p5_ASAP7_75t_R register___U5638 ( .A(register__net89877), .B(register__n1886), .Y(register__n2526) );
  OR2x2_ASAP7_75t_R register___U5639 ( .A(register__net93375), .B(register__n1683), .Y(register__n2306) );
  NOR2x1p5_ASAP7_75t_R register___U5640 ( .A(register__net104679), .B(register__n2490), .Y(register__n2491) );
  AND2x2_ASAP7_75t_R register___U5641 ( .A(register__n4444), .B(register__n2779), .Y(register__n2746) );
  OA211x2_ASAP7_75t_R register___U5642 ( .A1(register__C6423_net60749), .A2(register__n713), .B(register__n2512), .C(
        n2514), .Y(register__n2513) );
  INVx2_ASAP7_75t_R register___U5643 ( .A(register__n2513), .Y(register__n1891) );
  HB1xp67_ASAP7_75t_R register___U5644 ( .A(register__n2672), .Y(register__n1892) );
  NOR2xp67_ASAP7_75t_R register___U5645 ( .A(register__n2730), .B(register__n2702), .Y(register__n2733) );
  AO221x2_ASAP7_75t_R register___U5646 ( .A1(register__n233), .A2(register__net89997), .B1(register__n1226), .B2(
        net93741), .C(register__n2392), .Y(register__n2409) );
  INVx1_ASAP7_75t_R register___U5647 ( .A(register__n2409), .Y(register__n1893) );
  INVxp33_ASAP7_75t_R register___U5648 ( .A(register__n2026), .Y(register__n1894) );
  HB1xp67_ASAP7_75t_R register___U5649 ( .A(register__n1998), .Y(register__n1895) );
  HB1xp67_ASAP7_75t_R register___U5650 ( .A(register__n2562), .Y(register__n1896) );
  OA22x2_ASAP7_75t_R register___U5651 ( .A1(register__net150042), .A2(register__n2700), .B1(register__n2699), .B2(
        n_cell_124679_net155985), .Y(register__n2727) );
  INVx2_ASAP7_75t_R register___U5652 ( .A(register__n2727), .Y(register__n1897) );
  HB1xp67_ASAP7_75t_R register___U5653 ( .A(register__net150887), .Y(register__n1898) );
  OA21x2_ASAP7_75t_R register___U5654 ( .A1(register__n2026), .A2(register__n2427), .B(register__n2447), .Y(register__n2446) );
  INVx3_ASAP7_75t_R register___U5655 ( .A(register__n2446), .Y(register__n1899) );
  INVx1_ASAP7_75t_R register___U5656 ( .A(register__n2398), .Y(register__n1900) );
  OA221x2_ASAP7_75t_R register___U5657 ( .A1(register__C6422_net59965), .A2(register__n1800), .B1(
        C6423_net60880), .B2(register__n1114), .C(register__n2719), .Y(register__n2720) );
  INVx1_ASAP7_75t_R register___U5658 ( .A(register__n2720), .Y(register__n1902) );
  INVxp33_ASAP7_75t_R register___U5659 ( .A(register__n2075), .Y(register__n11571) );
  INVx1_ASAP7_75t_R register___U5660 ( .A(register__n6111), .Y(register__n2124) );
  INVx2_ASAP7_75t_R register___U5661 ( .A(register__n12072), .Y(register__n12052) );
  INVx1_ASAP7_75t_R register___U5662 ( .A(register__n9987), .Y(register__n2077) );
  INVx1_ASAP7_75t_R register___U5663 ( .A(register__n8765), .Y(register__n2076) );
  INVx1_ASAP7_75t_R register___U5664 ( .A(register__n9931), .Y(register__n2214) );
  INVx1_ASAP7_75t_R register___U5665 ( .A(register__n10471), .Y(register__n2199) );
  INVx1_ASAP7_75t_R register___U5666 ( .A(register__n9323), .Y(register__n2091) );
  INVx1_ASAP7_75t_R register___U5667 ( .A(register__n9915), .Y(register__n2126) );
  NOR4xp25_ASAP7_75t_R register___U5668 ( .A(register__n2722), .B(register__n2692), .C(register__n2725), .D(register__n2728), .Y(
        n2729) );
  INVx1_ASAP7_75t_R register___U5669 ( .A(register__n6892), .Y(register__n2090) );
  INVx1_ASAP7_75t_R register___U5670 ( .A(register__n8105), .Y(register__n2123) );
  INVx1_ASAP7_75t_R register___U5671 ( .A(register__n13326), .Y(register__n2039) );
  INVx1_ASAP7_75t_R register___U5672 ( .A(register__n13345), .Y(register__n2065) );
  INVx1_ASAP7_75t_R register___U5673 ( .A(register__n13138), .Y(register__n2055) );
  INVx1_ASAP7_75t_R register___U5674 ( .A(register__n13022), .Y(register__n2070) );
  INVx1_ASAP7_75t_R register___U5675 ( .A(register__n13114), .Y(register__n2036) );
  INVx1_ASAP7_75t_R register___U5676 ( .A(register__n13172), .Y(register__n2050) );
  INVx1_ASAP7_75t_R register___U5677 ( .A(register__n12651), .Y(register__n2054) );
  INVx1_ASAP7_75t_R register___U5678 ( .A(register__n13374), .Y(register__n2069) );
  INVx1_ASAP7_75t_R register___U5679 ( .A(register__n12910), .Y(register__n2051) );
  INVx1_ASAP7_75t_R register___U5680 ( .A(register__n12648), .Y(register__n2030) );
  INVx1_ASAP7_75t_R register___U5681 ( .A(register__n13338), .Y(register__n2044) );
  INVx1_ASAP7_75t_R register___U5682 ( .A(register__n13348), .Y(register__n2047) );
  INVx1_ASAP7_75t_R register___U5683 ( .A(register__n13357), .Y(register__n2057) );
  INVx1_ASAP7_75t_R register___U5684 ( .A(register__n12761), .Y(register__n2048) );
  INVx1_ASAP7_75t_R register___U5685 ( .A(register__n13186), .Y(register__n2027) );
  INVx1_ASAP7_75t_R register___U5686 ( .A(register__n13362), .Y(register__n2074) );
  INVx1_ASAP7_75t_R register___U5687 ( .A(register__n13343), .Y(register__n2067) );
  INVx1_ASAP7_75t_R register___U5688 ( .A(register__n13185), .Y(register__n2029) );
  INVx1_ASAP7_75t_R register___U5689 ( .A(register__n12699), .Y(register__n2046) );
  INVx1_ASAP7_75t_R register___U5690 ( .A(register__n12986), .Y(register__n2031) );
  INVx1_ASAP7_75t_R register___U5691 ( .A(register__n12700), .Y(register__n2034) );
  INVx1_ASAP7_75t_R register___U5692 ( .A(register__n13314), .Y(register__n2043) );
  INVx1_ASAP7_75t_R register___U5693 ( .A(register__n12955), .Y(register__n2032) );
  INVx1_ASAP7_75t_R register___U5694 ( .A(register__n13363), .Y(register__n2049) );
  INVx1_ASAP7_75t_R register___U5695 ( .A(register__n13356), .Y(register__n2063) );
  INVx1_ASAP7_75t_R register___U5696 ( .A(register__n13385), .Y(register__n2072) );
  INVx1_ASAP7_75t_R register___U5697 ( .A(register__n13280), .Y(register__n2033) );
  INVx1_ASAP7_75t_R register___U5698 ( .A(register__n13140), .Y(register__n2061) );
  INVx1_ASAP7_75t_R register___U5699 ( .A(register__n13382), .Y(register__n2062) );
  INVx1_ASAP7_75t_R register___U5700 ( .A(register__n12715), .Y(register__n2052) );
  INVx1_ASAP7_75t_R register___U5701 ( .A(register__n12916), .Y(register__n2059) );
  INVx1_ASAP7_75t_R register___U5702 ( .A(register__n13004), .Y(register__n2042) );
  INVx1_ASAP7_75t_R register___U5703 ( .A(register__n12694), .Y(register__n2058) );
  INVx1_ASAP7_75t_R register___U5704 ( .A(register__n12604), .Y(register__n2056) );
  INVx1_ASAP7_75t_R register___U5705 ( .A(register__n12592), .Y(register__n2040) );
  INVx1_ASAP7_75t_R register___U5706 ( .A(register__n12714), .Y(register__n2037) );
  INVx1_ASAP7_75t_R register___U5707 ( .A(register__n13372), .Y(register__n2073) );
  INVx1_ASAP7_75t_R register___U5708 ( .A(register__n13025), .Y(register__n2071) );
  INVx1_ASAP7_75t_R register___U5709 ( .A(register__n13359), .Y(register__n2035) );
  INVx1_ASAP7_75t_R register___U5710 ( .A(register__n12688), .Y(register__n2045) );
  NOR2x1_ASAP7_75t_R register___U5711 ( .A(register__n1907), .B(register__n1908), .Y(register__n13141) );
  NOR2x1_ASAP7_75t_R register___U5712 ( .A(register__n1266), .B(register__net64756), .Y(register__n1907) );
  NOR2x1_ASAP7_75t_R register___U5713 ( .A(register__n3335), .B(register__net90793), .Y(register__n1908) );
  INVx1_ASAP7_75t_R register___U5714 ( .A(register__n12913), .Y(register__n2041) );
  INVx1_ASAP7_75t_R register___U5715 ( .A(register__n13141), .Y(register__n2068) );
  BUFx12f_ASAP7_75t_R register___U5716 ( .A(register__net105921), .Y(register__net90793) );
  INVx1_ASAP7_75t_R register___U5717 ( .A(register__n13008), .Y(register__n2038) );
  INVx1_ASAP7_75t_R register___U5718 ( .A(register__n13344), .Y(register__n2066) );
  INVx1_ASAP7_75t_R register___U5719 ( .A(register__n13346), .Y(register__n2064) );
  INVx1_ASAP7_75t_R register___U5720 ( .A(register__n13277), .Y(register__n2060) );
  INVx2_ASAP7_75t_R register___U5721 ( .A(register__n1910), .Y(register__n1911) );
  INVxp33_ASAP7_75t_R register___U5722 ( .A(register__n1912), .Y(register__n1914) );
  INVxp67_ASAP7_75t_R register___U5723 ( .A(register__n2808), .Y(register__n1920) );
  INVxp33_ASAP7_75t_R register___U5724 ( .A(register__n1923), .Y(register__n1924) );
  INVxp33_ASAP7_75t_R register___U5725 ( .A(register__n1923), .Y(register__n1925) );
  HB1xp67_ASAP7_75t_R register___U5726 ( .A(register__n2803), .Y(register__n2810) );
  INVxp33_ASAP7_75t_R register___U5727 ( .A(register__n1927), .Y(register__n1928) );
  INVxp33_ASAP7_75t_R register___U5728 ( .A(register__n1927), .Y(register__n1929) );
  HB1xp67_ASAP7_75t_R register___U5729 ( .A(register__n2803), .Y(register__n2811) );
  INVxp33_ASAP7_75t_R register___U5730 ( .A(register__n1931), .Y(register__n1932) );
  INVxp33_ASAP7_75t_R register___U5731 ( .A(register__n1934), .Y(register__n1935) );
  INVxp33_ASAP7_75t_R register___U5732 ( .A(register__n1934), .Y(register__n1936) );
  INVxp33_ASAP7_75t_R register___U5733 ( .A(register__n1938), .Y(register__n1939) );
  INVxp33_ASAP7_75t_R register___U5734 ( .A(register__n1938), .Y(register__n1940) );
  INVxp33_ASAP7_75t_R register___U5735 ( .A(register__n1942), .Y(register__n1943) );
  INVxp33_ASAP7_75t_R register___U5736 ( .A(register__n1942), .Y(register__n1944) );
  HB1xp67_ASAP7_75t_R register___U5737 ( .A(register__n2804), .Y(register__n2815) );
  BUFx12f_ASAP7_75t_R register___U5738 ( .A(register__net117948), .Y(register__n1949) );
  INVx1_ASAP7_75t_R register___U5739 ( .A(register__net66316), .Y(register__n2462) );
  BUFx6f_ASAP7_75t_R register___U5740 ( .A(register__net66316), .Y(register__net66320) );
  INVx3_ASAP7_75t_R register___U5741 ( .A(register__n1949), .Y(register__n2185) );
  NAND2x1p5_ASAP7_75t_R register___U5742 ( .A(register__n2741), .B(register__n1990), .Y(register__n1955) );
  INVx2_ASAP7_75t_R register___U5743 ( .A(register__n10084), .Y(register__n2741) );
  BUFx6f_ASAP7_75t_R register___U5744 ( .A(register__n2021), .Y(register__n1990) );
  INVx2_ASAP7_75t_R register___U5745 ( .A(register__n1887), .Y(register__n2805) );
  BUFx6f_ASAP7_75t_R register___U5746 ( .A(register__n4894), .Y(register__n7059) );
  INVx3_ASAP7_75t_R register___U5747 ( .A(register__n7059), .Y(register__n1969) );
  INVx3_ASAP7_75t_R register___U5748 ( .A(register__n1969), .Y(register__n2206) );
  HB1xp67_ASAP7_75t_R register___U5749 ( .A(register__C6423_net61333), .Y(register__n2004) );
  NAND2xp5_ASAP7_75t_R register___U5750 ( .A(register__net90401), .B(register__net150051), .Y(register__n2502) );
  BUFx12f_ASAP7_75t_R register___U5751 ( .A(register__n11903), .Y(register__n11820) );
  INVxp33_ASAP7_75t_R register___U5752 ( .A(register__n2010), .Y(register__n2012) );
  OA22x2_ASAP7_75t_R register___U5753 ( .A1(register__n2076), .A2(register__C6423_net72243), .B1(register__n2077), .B2(
        n_cell_124679_net155985), .Y(register__n2075) );
  INVxp67_ASAP7_75t_R register___U5754 ( .A(register__n2897), .Y(register__n3999) );
  AO22x1_ASAP7_75t_R register___U5755 ( .A1(register__n9660), .A2(register__net122601), .B1(register__n9989), .B2(
        net125803), .Y(register__n11552) );
  AO22x1_ASAP7_75t_R register___U5756 ( .A1(register__n8528), .A2(register__net122601), .B1(register__n9433), .B2(
        net125803), .Y(register__n11377) );
  HB1xp67_ASAP7_75t_R register___U5757 ( .A(register__net122410), .Y(register__net122406) );
  INVxp67_ASAP7_75t_R register___U5758 ( .A(register__n3830), .Y(register__n6728) );
  INVxp67_ASAP7_75t_R register___U5759 ( .A(register__n4295), .Y(register__n7892) );
  HB1xp67_ASAP7_75t_R register___U5760 ( .A(register__n4296), .Y(register__n4295) );
  HB1xp67_ASAP7_75t_R register___U5761 ( .A(register__n5796), .Y(register__n5795) );
  INVxp67_ASAP7_75t_R register___U5762 ( .A(register__n3899), .Y(register__n6182) );
  HB1xp67_ASAP7_75t_R register___U5763 ( .A(register__n3900), .Y(register__n3899) );
  HB1xp67_ASAP7_75t_R register___U5764 ( .A(register__n11910), .Y(register__n3718) );
  HB1xp67_ASAP7_75t_R register___U5765 ( .A(register__n3718), .Y(register__n3717) );
  BUFx12f_ASAP7_75t_R register___U5766 ( .A(register__n7087), .Y(register__n3690) );
  BUFx6f_ASAP7_75t_R register___U5767 ( .A(register__n6464), .Y(register__n4037) );
  INVx1_ASAP7_75t_R register___U5768 ( .A(register__n12598), .Y(register__n2079) );
  HB1xp67_ASAP7_75t_R register___U5769 ( .A(register__n12934), .Y(register__n3965) );
  HB1xp67_ASAP7_75t_R register___U5770 ( .A(register__n3854), .Y(register__n3853) );
  HB1xp67_ASAP7_75t_R register___U5771 ( .A(register__n12590), .Y(register__n3854) );
  INVxp67_ASAP7_75t_R register___U5772 ( .A(register__n4785), .Y(register__n5374) );
  HB1xp67_ASAP7_75t_R register___U5773 ( .A(register__n4786), .Y(register__n4785) );
  AO22x1_ASAP7_75t_R register___U5774 ( .A1(register__n9863), .A2(register__net110414), .B1(register__n7229), .B2(
        net125797), .Y(register__n11362) );
  AO22x1_ASAP7_75t_R register___U5775 ( .A1(register__n9627), .A2(register__net110414), .B1(register__n10090), .B2(
        n1074), .Y(register__n11337) );
  HB1xp67_ASAP7_75t_R register___U5776 ( .A(register__n11536), .Y(register__n3055) );
  AO22x1_ASAP7_75t_R register___U5777 ( .A1(register__n9794), .A2(register__net110414), .B1(register__n10197), .B2(
        net117889), .Y(register__n11424) );
  NOR2xp33_ASAP7_75t_R register___U5778 ( .A(register__n9798), .B(register__n214), .Y(register__n2083) );
  INVxp67_ASAP7_75t_R register___U5779 ( .A(register__n12678), .Y(register__n2084) );
  INVx1_ASAP7_75t_R register___U5780 ( .A(register__n12600), .Y(register__n2085) );
  HB1xp67_ASAP7_75t_R register___U5781 ( .A(register__n13131), .Y(register__n2897) );
  HB1xp67_ASAP7_75t_R register___U5782 ( .A(register__n13165), .Y(register__n3967) );
  HB1xp67_ASAP7_75t_R register___U5783 ( .A(register__n10602), .Y(register__n2845) );
  INVxp67_ASAP7_75t_R register___U5784 ( .A(register__n2845), .Y(register__n3820) );
  HB1xp67_ASAP7_75t_R register___U5785 ( .A(register__n12582), .Y(register__n4786) );
  INVx1_ASAP7_75t_R register___U5786 ( .A(register__n11425), .Y(register__n2087) );
  AND2x2_ASAP7_75t_R register___U5787 ( .A(register__n2190), .B(register__n11406), .Y(register__n2088) );
  AND3x1_ASAP7_75t_R register___U5788 ( .A(register__n2088), .B(register__n11408), .C(register__n11407), .Y(register__n9154) );
  NOR3xp33_ASAP7_75t_R register___U5789 ( .A(register__n592), .B(register__n8340), .C(register__n8339), .Y(register__n2190) );
  HB1xp67_ASAP7_75t_R register___U5790 ( .A(register__n3831), .Y(register__n3830) );
  INVxp67_ASAP7_75t_R register___U5791 ( .A(register__n6795), .Y(register__n8677) );
  CKINVDCx10_ASAP7_75t_R register___U5792 ( .A(register__net63152), .Y(register__net97365) );
  CKINVDCx10_ASAP7_75t_R register___U5793 ( .A(register__net63186), .Y(register__net63152) );
  AND2x2_ASAP7_75t_R register___U5794 ( .A(register__n3440), .B(register__n6425), .Y(register__n2089) );
  AO22x1_ASAP7_75t_R register___U5795 ( .A1(register__n10499), .A2(register__net129017), .B1(register__n10454), .B2(
        n422), .Y(register__n11190) );
  INVxp33_ASAP7_75t_R register___U5796 ( .A(register__n11314), .Y(register__n5354) );
  INVx2_ASAP7_75t_R register___U5797 ( .A(register__n4812), .Y(register__n2203) );
  OAI22xp33_ASAP7_75t_R register___U5798 ( .A1(register__n2090), .A2(register__n793), .B1(register__n2091), .B2(
        net150880), .Y(register__n11444) );
  AND2x2_ASAP7_75t_R register___U5799 ( .A(register__n6549), .B(register__n5598), .Y(register__n2092) );
  INVxp33_ASAP7_75t_R register___U5800 ( .A(register__net66594), .Y(register__n2093) );
  INVxp33_ASAP7_75t_R register___U5801 ( .A(register__net73061), .Y(register__n2097) );
  INVx1_ASAP7_75t_R register___U5802 ( .A(register__net104558), .Y(register__n2103) );
  INVx1_ASAP7_75t_R register___U5803 ( .A(register__n2103), .Y(register__n2104) );
  INVx1_ASAP7_75t_R register___U5804 ( .A(register__n2107), .Y(register__n2108) );
  INVx2_ASAP7_75t_R register___U5805 ( .A(register__n2109), .Y(register__n2110) );
  INVx1_ASAP7_75t_R register___U5806 ( .A(register__n2113), .Y(register__n2114) );
  INVx2_ASAP7_75t_R register___U5807 ( .A(register__net104558), .Y(register__net73015) );
  HB1xp67_ASAP7_75t_R register___U5808 ( .A(register__net66594), .Y(register__net146710) );
  CKINVDCx10_ASAP7_75t_R register___U5809 ( .A(register__net141879), .Y(register__net73061) );
  INVx2_ASAP7_75t_R register___U5810 ( .A(register__net73015), .Y(register__net66582) );
  INVx4_ASAP7_75t_R register___U5811 ( .A(register__net73019), .Y(register__net66574) );
  HB1xp67_ASAP7_75t_R register___U5812 ( .A(register__n5435), .Y(register__n5434) );
  AO22x1_ASAP7_75t_R register___U5813 ( .A1(register__n9764), .A2(register__n481), .B1(register__n10257), .B2(register__n647), 
        .Y(register__n11599) );
  AO22x1_ASAP7_75t_R register___U5814 ( .A1(register__net88416), .A2(register__n481), .B1(register__net88504), .B2(
        C6423_net61348), .Y(register__n11616) );
  AO22x1_ASAP7_75t_R register___U5815 ( .A1(register__n9907), .A2(register__n481), .B1(register__n10210), .B2(register__n636), 
        .Y(register__n11427) );
  AO22x1_ASAP7_75t_R register___U5816 ( .A1(register__n9333), .A2(register__n482), .B1(register__n8789), .B2(register__n637), .Y(
        n11446) );
  INVxp67_ASAP7_75t_R register___U5817 ( .A(register__n6508), .Y(register__n7026) );
  BUFx12f_ASAP7_75t_R register___U5818 ( .A(register__net144981), .Y(register__net64446) );
  HB1xp67_ASAP7_75t_R register___U5819 ( .A(register__n11381), .Y(register__n5435) );
  INVxp33_ASAP7_75t_R register___U5820 ( .A(register__n5597), .Y(register__n6547) );
  INVxp67_ASAP7_75t_R register___U5821 ( .A(register__n12661), .Y(register__n7618) );
  INVxp33_ASAP7_75t_R register___U5822 ( .A(register__n4698), .Y(register__n7303) );
  HB1xp67_ASAP7_75t_R register___U5823 ( .A(register__n7303), .Y(register__n4700) );
  BUFx12f_ASAP7_75t_R register___U5824 ( .A(register__net128003), .Y(register__net136856) );
  HB1xp67_ASAP7_75t_R register___U5825 ( .A(register__n13044), .Y(register__n3831) );
  INVxp33_ASAP7_75t_R register___U5826 ( .A(register__n3238), .Y(register__n6424) );
  HB1xp67_ASAP7_75t_R register___U5827 ( .A(register__n6712), .Y(register__n4720) );
  HB1xp67_ASAP7_75t_R register___U5828 ( .A(register__n13096), .Y(register__n4085) );
  HB1xp67_ASAP7_75t_R register___U5829 ( .A(register__n12107), .Y(register__n12094) );
  INVxp33_ASAP7_75t_R register___U5830 ( .A(register__n4679), .Y(register__n7881) );
  HB1xp67_ASAP7_75t_R register___U5831 ( .A(register__n7881), .Y(register__n4681) );
  OAI22xp33_ASAP7_75t_R register___U5832 ( .A1(register__n2125), .A2(register__net150042), .B1(register__n2126), .B2(
        n2023), .Y(register__n11575) );
  CKINVDCx20_ASAP7_75t_R register___U5833 ( .A(register__n9668), .Y(register__n2125) );
  INVxp67_ASAP7_75t_R register___U5834 ( .A(register__n11122), .Y(register__n8747) );
  HB1xp67_ASAP7_75t_R register___U5835 ( .A(register__n4224), .Y(register__n4223) );
  HB1xp67_ASAP7_75t_R register___U5836 ( .A(register__n12662), .Y(register__n6796) );
  HB1xp67_ASAP7_75t_R register___U5837 ( .A(register__n6424), .Y(register__n3240) );
  INVx1_ASAP7_75t_R register___U5838 ( .A(register__n12732), .Y(register__n2128) );
  HB1xp67_ASAP7_75t_R register___U5839 ( .A(register__n11443), .Y(register__n4224) );
  HB1xp67_ASAP7_75t_R register___U5840 ( .A(register__n6796), .Y(register__n6795) );
  AO22x1_ASAP7_75t_R register___U5841 ( .A1(register__n9595), .A2(register__net121619), .B1(register__n10016), .B2(
        net126625), .Y(register__n10545) );
  AO22x1_ASAP7_75t_R register___U5842 ( .A1(register__n7800), .A2(register__n1771), .B1(register__n8133), .B2(register__net126625), .Y(register__n10653) );
  HB1xp67_ASAP7_75t_R register___U5843 ( .A(register__n6509), .Y(register__n6508) );
  INVxp33_ASAP7_75t_R register___U5844 ( .A(register__n4096), .Y(register__n8580) );
  CKINVDCx10_ASAP7_75t_R register___U5845 ( .A(register__net63154), .Y(register__net91738) );
  AO22x1_ASAP7_75t_R register___U5846 ( .A1(register__n9280), .A2(register__net122579), .B1(register__n9933), .B2(register__n1895), .Y(register__n11491) );
  AO22x1_ASAP7_75t_R register___U5847 ( .A1(register__n8194), .A2(register__n1966), .B1(register__n10233), .B2(register__n767), 
        .Y(register__n11381) );
  HB1xp67_ASAP7_75t_R register___U5848 ( .A(register__n5919), .Y(register__n5436) );
  INVxp67_ASAP7_75t_R register___U5849 ( .A(register__n4016), .Y(register__n6407) );
  OAI22xp33_ASAP7_75t_R register___U5850 ( .A1(register__n2130), .A2(register__net150046), .B1(register__n2131), .B2(
        n2023), .Y(register__n11633) );
  CKINVDCx20_ASAP7_75t_R register___U5851 ( .A(register__n9867), .Y(register__n2130) );
  CKINVDCx20_ASAP7_75t_R register___U5852 ( .A(register__n10291), .Y(register__n2131) );
  NOR2xp67_ASAP7_75t_R register___U5853 ( .A(register__net99861), .B(register__n2701), .Y(register__n2702) );
  AO22x1_ASAP7_75t_R register___U5854 ( .A1(register__n9335), .A2(register__net98137), .B1(register__n9355), .B2(register__n767), 
        .Y(register__n11443) );
  HB1xp67_ASAP7_75t_R register___U5855 ( .A(register__n11467), .Y(register__n5597) );
  INVxp67_ASAP7_75t_R register___U5856 ( .A(register__n5035), .Y(register__n2132) );
  HB1xp67_ASAP7_75t_R register___U5857 ( .A(register__n12109), .Y(register__n5035) );
  INVxp33_ASAP7_75t_R register___U5858 ( .A(register__n3052), .Y(register__n7879) );
  HB1xp67_ASAP7_75t_R register___U5859 ( .A(register__n12650), .Y(register__n6509) );
  INVxp33_ASAP7_75t_R register___U5860 ( .A(register__net66614), .Y(register__net66594) );
  INVx6_ASAP7_75t_R register___U5861 ( .A(register__n3502), .Y(register__n12082) );
  BUFx12f_ASAP7_75t_R register___U5862 ( .A(register__n3362), .Y(register__n3502) );
  INVx1_ASAP7_75t_R register___U5863 ( .A(register__n13229), .Y(register__n2133) );
  HB1xp67_ASAP7_75t_R register___U5864 ( .A(register__n6547), .Y(register__n5598) );
  HB1xp67_ASAP7_75t_R register___U5865 ( .A(register__n3975), .Y(register__n3974) );
  INVxp67_ASAP7_75t_R register___U5866 ( .A(register__n3974), .Y(register__n6187) );
  INVxp67_ASAP7_75t_R register___U5867 ( .A(register__n4297), .Y(register__n7032) );
  HB1xp67_ASAP7_75t_R register___U5868 ( .A(register__n13261), .Y(register__n4297) );
  HB1xp67_ASAP7_75t_R register___U5869 ( .A(register__n5354), .Y(register__n3919) );
  HB1xp67_ASAP7_75t_R register___U5870 ( .A(register__n4699), .Y(register__n4698) );
  HB1xp67_ASAP7_75t_R register___U5871 ( .A(register__n11401), .Y(register__n4699) );
  BUFx2_ASAP7_75t_R register___U5872 ( .A(register__n4262), .Y(register__n4261) );
  HB1xp67_ASAP7_75t_R register___U5873 ( .A(register__n4680), .Y(register__n4679) );
  AO22x1_ASAP7_75t_R register___U5874 ( .A1(register__n9260), .A2(register__C6423_net61333), .B1(register__n9923), .B2(
        n767), .Y(register__n11255) );
  HB1xp67_ASAP7_75t_R register___U5875 ( .A(register__n11792), .Y(register__n11788) );
  HB1xp67_ASAP7_75t_R register___U5876 ( .A(register__n11792), .Y(register__n11793) );
  BUFx12f_ASAP7_75t_R register___U5877 ( .A(register__n11785), .Y(register__n11787) );
  HB1xp67_ASAP7_75t_R register___U5878 ( .A(register__n11794), .Y(register__n11786) );
  HB1xp67_ASAP7_75t_R register___U5879 ( .A(register__n11798), .Y(register__n11784) );
  HB1xp67_ASAP7_75t_R register___U5880 ( .A(register__n4017), .Y(register__n4016) );
  HB1xp67_ASAP7_75t_R register___U5881 ( .A(register__n11489), .Y(register__n4017) );
  INVxp67_ASAP7_75t_R register___U5882 ( .A(register__n4823), .Y(register__n6431) );
  AO22x1_ASAP7_75t_R register___U5883 ( .A1(register__n9883), .A2(register__n1966), .B1(register__n10317), .B2(register__n767), 
        .Y(register__n11467) );
  AOI21xp33_ASAP7_75t_R register___U5884 ( .A1(register__net128096), .A2(register__net93753), .B(register__n2631), .Y(
        n2628) );
  AO22x1_ASAP7_75t_R register___U5885 ( .A1(register__n9282), .A2(register__n921), .B1(register__n10152), .B2(register__net150887), .Y(register__n11403) );
  AO22x1_ASAP7_75t_R register___U5886 ( .A1(register__n6621), .A2(register__n926), .B1(register__n9935), .B2(register__net150892), 
        .Y(register__n11338) );
  AO22x1_ASAP7_75t_R register___U5887 ( .A1(register__n9913), .A2(register__n932), .B1(register__n10216), .B2(register__n770), 
        .Y(register__n11697) );
  INVx6_ASAP7_75t_R register___U5888 ( .A(register__net138526), .Y(register__net120805) );
  AO22x1_ASAP7_75t_R register___U5889 ( .A1(register__n6981), .A2(register__n934), .B1(register__net150889), .B2(register__n10218), .Y(register__n11425) );
  HB1xp67_ASAP7_75t_R register___U5890 ( .A(register__net138612), .Y(register__n2137) );
  HB1xp67_ASAP7_75t_R register___U5891 ( .A(register__net138612), .Y(register__n2138) );
  HB1xp67_ASAP7_75t_R register___U5892 ( .A(register__n3053), .Y(register__n3052) );
  BUFx5_ASAP7_75t_R register___U5893 ( .A(register__n7257), .Y(register__n12097) );
  BUFx12_ASAP7_75t_R register___U5894 ( .A(register__n7257), .Y(register__n12095) );
  NOR2xp67_ASAP7_75t_R register___U5895 ( .A(register__net130031), .B(register__n2537), .Y(register__n2539) );
  INVxp67_ASAP7_75t_R register___U5896 ( .A(register__n4702), .Y(register__n7268) );
  HB1xp67_ASAP7_75t_R register___U5897 ( .A(register__n11633), .Y(register__n4262) );
  HB1xp67_ASAP7_75t_R register___U5898 ( .A(register__n12520), .Y(register__n4823) );
  HB1xp67_ASAP7_75t_R register___U5899 ( .A(register__n11273), .Y(register__n4680) );
  AO22x1_ASAP7_75t_R register___U5900 ( .A1(register__net90829), .A2(register__n1894), .B1(register__net90145), .B2(
        n767), .Y(register__n11273) );
  HB1xp67_ASAP7_75t_R register___U5901 ( .A(register__n4097), .Y(register__n4096) );
  HB1xp67_ASAP7_75t_R register___U5902 ( .A(register__n8580), .Y(register__n4098) );
  INVxp33_ASAP7_75t_R register___U5903 ( .A(register__net74029), .Y(register__n2143) );
  INVx2_ASAP7_75t_R register___U5904 ( .A(register__net106927), .Y(register__net73985) );
  INVx2_ASAP7_75t_R register___U5905 ( .A(register__n4657), .Y(register__n6435) );
  BUFx3_ASAP7_75t_R register___U5906 ( .A(register__n4658), .Y(register__n4657) );
  INVxp67_ASAP7_75t_R register___U5907 ( .A(register__n7363), .Y(register__n9236) );
  HB1xp67_ASAP7_75t_R register___U5908 ( .A(register__n12703), .Y(register__n3549) );
  HB1xp67_ASAP7_75t_R register___U5909 ( .A(register__n11505), .Y(register__n4030) );
  INVxp67_ASAP7_75t_R register___U5910 ( .A(register__n3548), .Y(register__n5234) );
  HB1xp67_ASAP7_75t_R register___U5911 ( .A(register__n3549), .Y(register__n3548) );
  HB1xp67_ASAP7_75t_R register___U5912 ( .A(register__n11575), .Y(register__n4097) );
  AO22x1_ASAP7_75t_R register___U5913 ( .A1(register__n9286), .A2(register__n922), .B1(register__n10169), .B2(register__net150873), .Y(register__n11363) );
  HB1xp67_ASAP7_75t_R register___U5914 ( .A(register__n11539), .Y(register__n3053) );
  AO22x1_ASAP7_75t_R register___U5915 ( .A1(register__n9644), .A2(register__net109849), .B1(register__n9971), .B2(register__n643), 
        .Y(register__n11539) );
  HB1xp67_ASAP7_75t_R register___U5916 ( .A(register__n7364), .Y(register__n7363) );
  HB1xp67_ASAP7_75t_R register___U5917 ( .A(register__n3610), .Y(register__n3609) );
  HB1xp67_ASAP7_75t_R register___U5918 ( .A(register__n12708), .Y(register__n5774) );
  HB1xp67_ASAP7_75t_R register___U5919 ( .A(register__n4703), .Y(register__n4702) );
  BUFx12_ASAP7_75t_R register___U5920 ( .A(register__n3565), .Y(register__n12077) );
  INVxp67_ASAP7_75t_R register___U5921 ( .A(register__n3332), .Y(register__n8622) );
  HB1xp67_ASAP7_75t_R register___U5922 ( .A(register__n7268), .Y(register__n4704) );
  BUFx12f_ASAP7_75t_R register___U5923 ( .A(register__net140685), .Y(register__net63186) );
  HB1xp67_ASAP7_75t_R register___U5924 ( .A(register__n11512), .Y(register__n4703) );
  AND2x2_ASAP7_75t_R register___U5925 ( .A(register__n10518), .B(register__n830), .Y(register__n4127) );
  HB1xp67_ASAP7_75t_R register___U5926 ( .A(register__n4127), .Y(register__n11848) );
  AO22x1_ASAP7_75t_R register___U5927 ( .A1(register__n9824), .A2(register__n85), .B1(register__n10235), .B2(register__n422), .Y(
        n11511) );
  HB1xp67_ASAP7_75t_R register___U5928 ( .A(register__n11850), .Y(register__n2155) );
  BUFx6f_ASAP7_75t_R register___U5929 ( .A(register__n4374), .Y(register__n2984) );
  HB1xp67_ASAP7_75t_R register___U5930 ( .A(register__n3390), .Y(register__n11849) );
  HB1xp67_ASAP7_75t_R register___U5931 ( .A(register__n13167), .Y(register__n3975) );
  AO22x1_ASAP7_75t_R register___U5932 ( .A1(register__n9303), .A2(register__n1966), .B1(register__n6948), .B2(
        C6423_net61331), .Y(register__n11512) );
  HB1xp67_ASAP7_75t_R register___U5933 ( .A(register__n11662), .Y(register__n7364) );
  BUFx3_ASAP7_75t_R register___U5934 ( .A(register__n5786), .Y(register__n5785) );
  CKINVDCx11_ASAP7_75t_R register___U5935 ( .A(register__n4004), .Y(register__n12081) );
  INVx1_ASAP7_75t_R register___U5936 ( .A(register__n2956), .Y(register__n4593) );
  HB1xp67_ASAP7_75t_R register___U5937 ( .A(register__n7879), .Y(register__n3054) );
  HB1xp67_ASAP7_75t_R register___U5938 ( .A(register__n13115), .Y(register__n5760) );
  AO22x1_ASAP7_75t_R register___U5939 ( .A1(register__n9272), .A2(register__C6423_net68948), .B1(register__n10237), 
        .B2(register__n2001), .Y(register__n11505) );
  AO22x1_ASAP7_75t_R register___U5940 ( .A1(register__n9788), .A2(register__n1853), .B1(register__n10104), .B2(
        net123857), .Y(register__n11114) );
  AO22x1_ASAP7_75t_R register___U5941 ( .A1(register__n9891), .A2(register__n1853), .B1(register__n9321), .B2(register__net123857), .Y(register__n11138) );
  AO22x1_ASAP7_75t_R register___U5942 ( .A1(register__n9696), .A2(register__net129747), .B1(register__n9967), .B2(
        C6422_net70296), .Y(register__n10540) );
  HB1xp67_ASAP7_75t_R register___U5943 ( .A(register__n4346), .Y(register__n4345) );
  INVxp67_ASAP7_75t_R register___U5944 ( .A(register__n4345), .Y(register__n7312) );
  HB1xp67_ASAP7_75t_R register___U5945 ( .A(register__n3862), .Y(register__n3861) );
  INVxp67_ASAP7_75t_R register___U5946 ( .A(register__n3861), .Y(register__n5532) );
  HB1xp67_ASAP7_75t_R register___U5947 ( .A(register__n12809), .Y(register__n3610) );
  HB1xp67_ASAP7_75t_R register___U5948 ( .A(register__n3196), .Y(register__n3195) );
  INVxp67_ASAP7_75t_R register___U5949 ( .A(register__n3195), .Y(register__n4388) );
  HB1xp67_ASAP7_75t_R register___U5950 ( .A(register__n13369), .Y(register__n3196) );
  HB1xp67_ASAP7_75t_R register___U5951 ( .A(register__n2829), .Y(register__n11794) );
  INVx1_ASAP7_75t_R register___U5952 ( .A(register__n10581), .Y(register__n2158) );
  HB1xp67_ASAP7_75t_R register___U5953 ( .A(register__n10987), .Y(register__n4346) );
  AO22x1_ASAP7_75t_R register___U5954 ( .A1(register__n9843), .A2(register__n1853), .B1(register__n10122), .B2(
        net123857), .Y(register__n10987) );
  HB1xp67_ASAP7_75t_R register___U5955 ( .A(register__n11006), .Y(register__n3862) );
  AO22x1_ASAP7_75t_R register___U5956 ( .A1(register__net90813), .A2(register__C6422_net60422), .B1(register__net90061), 
        .B2(register__net123857), .Y(register__n11006) );
  NOR3x1_ASAP7_75t_R register___U5957 ( .A(register__n10753), .B(register__n5030), .C(register__n5028), .Y(register__n2778) );
  NAND4xp75_ASAP7_75t_R register___U5958 ( .A(register__n8219), .B(register__n8220), .C(register__n8218), .D(register__n5260), 
        .Y(register__n2161) );
  HB1xp67_ASAP7_75t_R register___U5959 ( .A(register__n6786), .Y(register__n6785) );
  INVxp67_ASAP7_75t_R register___U5960 ( .A(register__n6785), .Y(register__n8620) );
  AO22x1_ASAP7_75t_R register___U5961 ( .A1(register__n10501), .A2(register__n768), .B1(register__n9246), .B2(register__n75), .Y(
        n11145) );
  BUFx6f_ASAP7_75t_R register___U5962 ( .A(register__n1951), .Y(register__n3710) );
  OAI22xp5_ASAP7_75t_R register___U5963 ( .A1(register__net62660), .A2(register__n11889), .B1(register__n9246), .B2(
        n12500), .Y(register__n2211) );
  INVx1_ASAP7_75t_R register___U5964 ( .A(register__n13370), .Y(register__n2164) );
  INVx1_ASAP7_75t_R register___U5965 ( .A(register__n13377), .Y(register__n2165) );
  AO22x1_ASAP7_75t_R register___U5966 ( .A1(register__n9244), .A2(register__n77), .B1(register__n10444), .B2(register__n75), .Y(
        n10609) );
  HB1xp67_ASAP7_75t_R register___U5967 ( .A(register__n3333), .Y(register__n3332) );
  AO22x1_ASAP7_75t_R register___U5968 ( .A1(register__n9349), .A2(register__C6422_net60422), .B1(register__n9367), .B2(
        net123857), .Y(register__n11071) );
  AO22x1_ASAP7_75t_R register___U5969 ( .A1(register__n9766), .A2(register__net129747), .B1(register__n10114), .B2(
        net123857), .Y(register__n11027) );
  AO22x1_ASAP7_75t_R register___U5970 ( .A1(register__n9694), .A2(register__net129747), .B1(register__n9965), .B2(
        net139537), .Y(register__n10581) );
  AO22x1_ASAP7_75t_R register___U5971 ( .A1(register__n9690), .A2(register__C6422_net60422), .B1(register__n9961), .B2(
        net123857), .Y(register__n10626) );
  AO22x1_ASAP7_75t_R register___U5972 ( .A1(register__n9692), .A2(register__net129746), .B1(register__n9963), .B2(
        net139537), .Y(register__n10606) );
  AO22x1_ASAP7_75t_R register___U5973 ( .A1(register__net90629), .A2(register__C6422_net60422), .B1(register__net89010), 
        .B2(register__net123857), .Y(register__n11090) );
  AO22x1_ASAP7_75t_R register___U5974 ( .A1(register__n9684), .A2(register__net129747), .B1(register__n9955), .B2(
        net123857), .Y(register__n10943) );
  AO22x1_ASAP7_75t_R register___U5975 ( .A1(register__n9847), .A2(register__net129747), .B1(register__n10167), .B2(
        net123857), .Y(register__n10690) );
  HB1xp67_ASAP7_75t_R register___U5976 ( .A(register__n10584), .Y(register__n4448) );
  AO22x1_ASAP7_75t_R register___U5977 ( .A1(register__n9632), .A2(register__C6422_net60445), .B1(register__n10068), 
        .B2(register__C6422_net60443), .Y(register__n10584) );
  AO22x1_ASAP7_75t_R register___U5978 ( .A1(register__n10509), .A2(register__n38), .B1(register__n10511), .B2(register__n369), 
        .Y(register__n10946) );
  HB1xp67_ASAP7_75t_R register___U5979 ( .A(register__n12737), .Y(register__n3776) );
  AO22x1_ASAP7_75t_R register___U5980 ( .A1(register__n9258), .A2(register__n1867), .B1(register__net96692), .B2(register__n9995), 
        .Y(register__n10604) );
  HB1xp67_ASAP7_75t_R register___U5981 ( .A(register__n10604), .Y(register__n3129) );
  NAND2x1p5_ASAP7_75t_R register___U5982 ( .A(register__n6705), .B(register__n7943), .Y(register__n2253) );
  OAI22xp33_ASAP7_75t_R register___U5983 ( .A1(register__net63242), .A2(register__n576), .B1(register__net103568), .B2(
        n586), .Y(register__n2168) );
  INVx1_ASAP7_75t_R register___U5984 ( .A(register__n12857), .Y(register__n2169) );
  INVx1_ASAP7_75t_R register___U5985 ( .A(register__n12853), .Y(register__n2170) );
  INVx3_ASAP7_75t_R register___U5986 ( .A(register__n7060), .Y(register__n2207) );
  INVx3_ASAP7_75t_R register___U5987 ( .A(register__n11531), .Y(register__n7060) );
  INVx1_ASAP7_75t_R register___U5988 ( .A(register__n12847), .Y(register__n2171) );
  INVx1_ASAP7_75t_R register___U5989 ( .A(register__n12858), .Y(register__n2172) );
  INVx1_ASAP7_75t_R register___U5990 ( .A(register__n12848), .Y(register__n2173) );
  INVx1_ASAP7_75t_R register___U5991 ( .A(register__n12577), .Y(register__n2174) );
  INVx1_ASAP7_75t_R register___U5992 ( .A(register__n12562), .Y(register__n2175) );
  INVx1_ASAP7_75t_R register___U5993 ( .A(register__n12718), .Y(register__n2176) );
  HB1xp67_ASAP7_75t_R register___U5994 ( .A(register__n13177), .Y(register__n6259) );
  HB1xp67_ASAP7_75t_R register___U5995 ( .A(register__n4739), .Y(register__n4738) );
  INVx1_ASAP7_75t_R register___U5996 ( .A(register__n12781), .Y(register__n2177) );
  INVx1_ASAP7_75t_R register___U5997 ( .A(register__n12780), .Y(register__n2178) );
  INVx1_ASAP7_75t_R register___U5998 ( .A(register__n12785), .Y(register__n2179) );
  INVx1_ASAP7_75t_R register___U5999 ( .A(register__n12783), .Y(register__n2180) );
  INVx1_ASAP7_75t_R register___U6000 ( .A(register__n12790), .Y(register__n2181) );
  INVx1_ASAP7_75t_R register___U6001 ( .A(register__n12782), .Y(register__n2182) );
  INVx1_ASAP7_75t_R register___U6002 ( .A(register__n12777), .Y(register__n2183) );
  INVx1_ASAP7_75t_R register___U6003 ( .A(register__n12784), .Y(register__n2184) );
  NAND3x1_ASAP7_75t_R register___U6004 ( .A(register__n2784), .B(register__n11640), .C(register__n259), .Y(register__n2186) );
  OR2x2_ASAP7_75t_R register___U6005 ( .A(register__net139024), .B(register__n1687), .Y(register__n2189) );
  HB1xp67_ASAP7_75t_R register___U6006 ( .A(register__n11628), .Y(register__n4739) );
  HB1xp67_ASAP7_75t_R register___U6007 ( .A(register__n4203), .Y(register__n4202) );
  INVx1_ASAP7_75t_R register___U6008 ( .A(register__n13037), .Y(register__n2191) );
  INVx1_ASAP7_75t_R register___U6009 ( .A(register__n13031), .Y(register__n2192) );
  INVx1_ASAP7_75t_R register___U6010 ( .A(register__n13027), .Y(register__n2193) );
  INVx1_ASAP7_75t_R register___U6011 ( .A(register__n12854), .Y(register__n2194) );
  INVx1_ASAP7_75t_R register___U6012 ( .A(register__n11681), .Y(register__n2195) );
  AO22x1_ASAP7_75t_R register___U6013 ( .A1(register__n12271), .A2(register__n535), .B1(register__n2197), .B2(register__n1098), 
        .Y(register__n2196) );
  CKINVDCx20_ASAP7_75t_R register___U6014 ( .A(register__n9933), .Y(register__n2197) );
  NOR2xp67_ASAP7_75t_R register___U6015 ( .A(register__n2525), .B(register__n2526), .Y(register__C6423_net60964) );
  BUFx2_ASAP7_75t_R register___U6016 ( .A(register__net122897), .Y(register__net122896) );
  AO22x1_ASAP7_75t_R register___U6017 ( .A1(register__n12304), .A2(register__n3217), .B1(register__n2199), .B2(register__n2220), 
        .Y(register__n2198) );
  INVx1_ASAP7_75t_R register___U6018 ( .A(register__n13021), .Y(register__n2200) );
  AO22x1_ASAP7_75t_R register___U6019 ( .A1(register__n12359), .A2(register__n3605), .B1(register__n2202), .B2(register__n2220), 
        .Y(register__n2201) );
  CKINVDCx20_ASAP7_75t_R register___U6020 ( .A(register__n9382), .Y(register__n2202) );
  HB1xp67_ASAP7_75t_R register___U6021 ( .A(register__n13241), .Y(register__n6786) );
  NOR4xp75_ASAP7_75t_R register___U6022 ( .A(register__n7305), .B(register__n4813), .C(register__n4997), .D(register__n2203), .Y(
        n11035) );
  INVx1_ASAP7_75t_R register___U6023 ( .A(register__n10644), .Y(register__n2205) );
  INVx2_ASAP7_75t_R register___U6024 ( .A(register__n4725), .Y(register__n7935) );
  NOR4xp75_ASAP7_75t_R register___U6025 ( .A(register__n2206), .B(register__n4896), .C(register__n5309), .D(register__n2207), .Y(
        n11519) );
  INVx1_ASAP7_75t_R register___U6026 ( .A(register__n12832), .Y(register__n2208) );
  INVx1_ASAP7_75t_R register___U6027 ( .A(register__n12616), .Y(register__n2209) );
  INVx1_ASAP7_75t_R register___U6028 ( .A(register__n12612), .Y(register__n2210) );
  INVx1_ASAP7_75t_R register___U6029 ( .A(register__n11387), .Y(register__n2212) );
  BUFx3_ASAP7_75t_R register___U6030 ( .A(register__n11433), .Y(register__n5120) );
  AO22x1_ASAP7_75t_R register___U6031 ( .A1(register__n12332), .A2(register__n3306), .B1(register__n2214), .B2(register__n2220), 
        .Y(register__n2213) );
  INVx2_ASAP7_75t_R register___U6032 ( .A(register__n12332), .Y(register__n12319) );
  INVx1_ASAP7_75t_R register___U6033 ( .A(register__n10730), .Y(register__n2215) );
  NAND2xp67_ASAP7_75t_R register___U6034 ( .A(register__n8236), .B(register__n2789), .Y(register__n2217) );
  INVx1_ASAP7_75t_R register___U6035 ( .A(register__n12608), .Y(register__n2218) );
  BUFx3_ASAP7_75t_R register___U6036 ( .A(register__n11411), .Y(register__n5821) );
  INVx1_ASAP7_75t_R register___U6037 ( .A(register__n13028), .Y(register__n2221) );
  HB1xp67_ASAP7_75t_R register___U6038 ( .A(register__n12578), .Y(register__n4203) );
  INVx2_ASAP7_75t_R register___U6039 ( .A(register__n5296), .Y(register__n7607) );
  INVx1_ASAP7_75t_R register___U6040 ( .A(register__n12611), .Y(register__n2223) );
  BUFx3_ASAP7_75t_R register___U6041 ( .A(register__n11390), .Y(register__n5814) );
  INVx1_ASAP7_75t_R register___U6042 ( .A(register__n10985), .Y(register__n2224) );
  AO22x1_ASAP7_75t_R register___U6043 ( .A1(register__n9415), .A2(register__net104772), .B1(register__n7216), .B2(register__n1357), .Y(register__n10985) );
  AO22x1_ASAP7_75t_R register___U6044 ( .A1(register__net110090), .A2(register__n168), .B1(register__net89597), .B2(
        net108158), .Y(register__n10730) );
  AO22x1_ASAP7_75t_R register___U6045 ( .A1(register__n9786), .A2(register__net146144), .B1(register__n10185), .B2(
        net126602), .Y(register__n10644) );
  INVx2_ASAP7_75t_R register___U6046 ( .A(register__n8638), .Y(register__n2281) );
  INVx1_ASAP7_75t_R register___U6047 ( .A(register__n11134), .Y(register__n2225) );
  INVx1_ASAP7_75t_R register___U6048 ( .A(register__n13107), .Y(register__n2226) );
  INVx1_ASAP7_75t_R register___U6049 ( .A(register__C6423_net72243), .Y(register__C6423_net72253) );
  AND3x1_ASAP7_75t_R register___U6050 ( .A(register__n7002), .B(register__n7001), .C(register__n7000), .Y(register__n2790) );
  INVx2_ASAP7_75t_R register___U6051 ( .A(register__n5585), .Y(register__n7001) );
  AO22x1_ASAP7_75t_R register___U6052 ( .A1(register__n7438), .A2(register__n413), .B1(register__n6563), .B2(register__net126602), 
        .Y(register__n10872) );
  AND3x1_ASAP7_75t_R register___U6053 ( .A(register__n8217), .B(register__n22), .C(register__register__n2215), .Y(register__n2789) );
  INVxp67_ASAP7_75t_R register___U6054 ( .A(register__n12710), .Y(register__n2227) );
  INVx1_ASAP7_75t_R register___U6055 ( .A(register__n11347), .Y(register__n2228) );
  INVx1_ASAP7_75t_R register___U6056 ( .A(register__n12786), .Y(register__n2229) );
  INVx1_ASAP7_75t_R register___U6057 ( .A(register__n12792), .Y(register__n2230) );
  INVx1_ASAP7_75t_R register___U6058 ( .A(register__n12791), .Y(register__n2231) );
  INVxp33_ASAP7_75t_R register___U6059 ( .A(register__n5586), .Y(register__n7928) );
  NOR2xp67_ASAP7_75t_R register___U6060 ( .A(register__n2793), .B(register__n2794), .Y(register__n12710) );
  INVx1_ASAP7_75t_R register___U6061 ( .A(register__n12606), .Y(register__n2232) );
  HB1xp67_ASAP7_75t_R register___U6062 ( .A(register__n13234), .Y(register__n3582) );
  HB1xp67_ASAP7_75t_R register___U6063 ( .A(register__n13204), .Y(register__n5969) );
  INVx1_ASAP7_75t_R register___U6064 ( .A(register__n13020), .Y(register__n2236) );
  INVx1_ASAP7_75t_R register___U6065 ( .A(register__n13032), .Y(register__n2237) );
  HB1xp67_ASAP7_75t_R register___U6066 ( .A(register__n5587), .Y(register__n5586) );
  INVx1_ASAP7_75t_R register___U6067 ( .A(register__n12635), .Y(register__n2238) );
  INVx1_ASAP7_75t_R register___U6068 ( .A(register__n13013), .Y(register__n2239) );
  INVx1_ASAP7_75t_R register___U6069 ( .A(register__n13035), .Y(register__n2240) );
  INVx1_ASAP7_75t_R register___U6070 ( .A(register__n13030), .Y(register__n2241) );
  AO22x1_ASAP7_75t_R register___U6071 ( .A1(register__n7550), .A2(register__n39), .B1(register__n7842), .B2(
        C6422_net60399), .Y(register__n11134) );
  NOR2xp67_ASAP7_75t_R register___U6072 ( .A(register__n2759), .B(register__n2760), .Y(register__n13195) );
  NOR2x2_ASAP7_75t_R register___U6073 ( .A(register__n12145), .B(register__n978), .Y(register__n2759) );
  INVx1_ASAP7_75t_R register___U6074 ( .A(register__n13033), .Y(register__n2242) );
  INVx1_ASAP7_75t_R register___U6075 ( .A(register__n13225), .Y(register__n2243) );
  INVx1_ASAP7_75t_R register___U6076 ( .A(register__n12624), .Y(register__n2247) );
  INVx1_ASAP7_75t_R register___U6077 ( .A(register__n13251), .Y(register__n2248) );
  BUFx3_ASAP7_75t_R register___U6078 ( .A(register__n11684), .Y(register__n5477) );
  BUFx12f_ASAP7_75t_R register___U6079 ( .A(register__n12077), .Y(register__n12068) );
  INVx2_ASAP7_75t_R register___U6080 ( .A(register__n3012), .Y(register__n6196) );
  HB1xp67_ASAP7_75t_R register___U6081 ( .A(register__n11430), .Y(register__n8271) );
  AO22x1_ASAP7_75t_R register___U6082 ( .A1(register__n10491), .A2(register__net146144), .B1(register__n8785), .B2(
        net126601), .Y(register__n10667) );
  BUFx6f_ASAP7_75t_R register___U6083 ( .A(register__net104773), .Y(register__net104772) );
  NOR2x1p5_ASAP7_75t_R register___U6084 ( .A(register__n12060), .B(register__n339), .Y(register__n2780) );
  AO22x1_ASAP7_75t_R register___U6085 ( .A1(register__n9903), .A2(register__n1867), .B1(register__n10206), .B2(register__n1360), 
        .Y(register__n11112) );
  AO22x1_ASAP7_75t_R register___U6086 ( .A1(register__n10495), .A2(register__net91683), .B1(register__n1347), .B2(
        n10450), .Y(register__n10560) );
  AO22x1_ASAP7_75t_R register___U6087 ( .A1(register__net101003), .A2(register__net91683), .B1(register__net112298), 
        .B2(register__net96692), .Y(register__n10707) );
  AO22x1_ASAP7_75t_R register___U6088 ( .A1(register__n9411), .A2(register__n1867), .B1(register__n9997), .B2(register__net96692), 
        .Y(register__n10538) );
  BUFx3_ASAP7_75t_R register___U6089 ( .A(register__n13134), .Y(register__n2957) );
  INVx1_ASAP7_75t_R register___U6090 ( .A(register__n11508), .Y(register__n2251) );
  AO22x1_ASAP7_75t_R register___U6091 ( .A1(register__n9760), .A2(register__C6423_net72253), .B1(register__n10245), 
        .B2(register__net139058), .Y(register__n11508) );
  HB1xp67_ASAP7_75t_R register___U6092 ( .A(register__n13135), .Y(register__n3047) );
  HB1xp67_ASAP7_75t_R register___U6093 ( .A(register__n13145), .Y(register__n2942) );
  BUFx3_ASAP7_75t_R register___U6094 ( .A(register__n2957), .Y(register__n2956) );
  INVx1_ASAP7_75t_R register___U6095 ( .A(register__n11649), .Y(register__n2252) );
  AO22x1_ASAP7_75t_R register___U6096 ( .A1(register__n8811), .A2(register__net138603), .B1(register__n8819), .B2(
        net125803), .Y(register__n11649) );
  HB1xp67_ASAP7_75t_R register___U6097 ( .A(register__n12587), .Y(register__n3459) );
  HB1xp67_ASAP7_75t_R register___U6098 ( .A(register__n2843), .Y(register__n11792) );
  HB1xp67_ASAP7_75t_R register___U6099 ( .A(register__n13183), .Y(register__n5766) );
  INVxp33_ASAP7_75t_R register___U6100 ( .A(register__n4551), .Y(register__n8260) );
  INVx1_ASAP7_75t_R register___U6101 ( .A(register__n12609), .Y(register__n2255) );
  INVx1_ASAP7_75t_R register___U6102 ( .A(register__n12610), .Y(register__n2256) );
  HB1xp67_ASAP7_75t_R register___U6103 ( .A(register__n11798), .Y(register__n11789) );
  HB1xp67_ASAP7_75t_R register___U6104 ( .A(register__n11571), .Y(register__n4551) );
  INVx1_ASAP7_75t_R register___U6105 ( .A(register__n13052), .Y(register__n2257) );
  XNOR2xp5_ASAP7_75t_R register___U6106 ( .A(register__n410), .B(register__n5523), .Y(register__n12507) );
  BUFx3_ASAP7_75t_R register___U6107 ( .A(register__n7316), .Y(register__n4256) );
  BUFx3_ASAP7_75t_R register___U6108 ( .A(register__n8276), .Y(register__n5618) );
  HB1xp67_ASAP7_75t_R register___U6109 ( .A(register__n12902), .Y(register__n3272) );
  INVx1_ASAP7_75t_R register___U6110 ( .A(register__n11165), .Y(register__n2258) );
  INVx1_ASAP7_75t_R register___U6111 ( .A(register__n11629), .Y(register__n2259) );
  AO22x1_ASAP7_75t_R register___U6112 ( .A1(register__n9111), .A2(register__net137440), .B1(register__n10283), .B2(
        C6423_net68764), .Y(register__n11629) );
  HB1xp67_ASAP7_75t_R register___U6113 ( .A(register__n12990), .Y(register__n5269) );
  INVx1_ASAP7_75t_R register___U6114 ( .A(register__n13231), .Y(register__n2260) );
  NOR3x1_ASAP7_75t_R register___U6115 ( .A(register__n11659), .B(register__n2261), .C(register__n2262), .Y(register__n3721) );
  INVxp67_ASAP7_75t_R register___U6116 ( .A(register__n3109), .Y(register__n7652) );
  HB1xp67_ASAP7_75t_R register___U6117 ( .A(register__n3239), .Y(register__n3238) );
  INVx1_ASAP7_75t_R register___U6118 ( .A(register__n13125), .Y(register__n2263) );
  INVx1_ASAP7_75t_R register___U6119 ( .A(register__n13126), .Y(register__n2264) );
  INVx1_ASAP7_75t_R register___U6120 ( .A(register__n13127), .Y(register__n2265) );
  INVx1_ASAP7_75t_R register___U6121 ( .A(register__n13232), .Y(register__n2266) );
  HB1xp67_ASAP7_75t_R register___U6122 ( .A(register__n3110), .Y(register__n3109) );
  INVx1_ASAP7_75t_R register___U6123 ( .A(register__n12921), .Y(register__n2267) );
  INVx1_ASAP7_75t_R register___U6124 ( .A(register__n12944), .Y(register__n2268) );
  INVx1_ASAP7_75t_R register___U6125 ( .A(register__n12941), .Y(register__n2269) );
  INVxp67_ASAP7_75t_R register___U6126 ( .A(register__n12684), .Y(register__n2270) );
  INVx1_ASAP7_75t_R register___U6127 ( .A(register__n12675), .Y(register__n2273) );
  HB1xp67_ASAP7_75t_R register___U6128 ( .A(register__n13075), .Y(register__n4296) );
  HB1xp67_ASAP7_75t_R register___U6129 ( .A(register__n13099), .Y(register__n5796) );
  HB1xp67_ASAP7_75t_R register___U6130 ( .A(register__n12994), .Y(register__n3888) );
  INVxp67_ASAP7_75t_R register___U6131 ( .A(register__n3888), .Y(register__n6180) );
  HB1xp67_ASAP7_75t_R register___U6132 ( .A(register__n13222), .Y(register__n3900) );
  NOR2xp67_ASAP7_75t_R register___U6133 ( .A(register__n2786), .B(register__n2787), .Y(register__n12684) );
  NOR2x1p5_ASAP7_75t_R register___U6134 ( .A(register__n12061), .B(register__n197), .Y(register__n2786) );
  HB1xp67_ASAP7_75t_R register___U6135 ( .A(register__n4153), .Y(register__n4152) );
  INVxp67_ASAP7_75t_R register___U6136 ( .A(register__n4152), .Y(register__n6130) );
  INVxp67_ASAP7_75t_R register___U6137 ( .A(register__n13353), .Y(register__n7616) );
  HB1xp67_ASAP7_75t_R register___U6138 ( .A(register__n12977), .Y(register__n2922) );
  NOR3x1_ASAP7_75t_R register___U6139 ( .A(register__n2282), .B(register__n5157), .C(register__n2281), .Y(register__n2755) );
  AND2x2_ASAP7_75t_R register___U6140 ( .A(IF_ID_rs1[0]), .B(IF_ID_rs1[1]), 
        .Y(register__n11136) );
  INVx1_ASAP7_75t_R register___U6141 ( .A(register__n10570), .Y(register__n9186) );
  INVx1_ASAP7_75t_R register___U6142 ( .A(register__n13228), .Y(register__n2283) );
  INVx1_ASAP7_75t_R register___U6143 ( .A(register__n13227), .Y(register__n2284) );
  HB1xp67_ASAP7_75t_R register___U6144 ( .A(register__n13339), .Y(register__n3898) );
  HB1xp67_ASAP7_75t_R register___U6145 ( .A(register__n13352), .Y(register__n4153) );
  INVx1_ASAP7_75t_R register___U6146 ( .A(register__n13337), .Y(register__n2287) );
  INVx1_ASAP7_75t_R register___U6147 ( .A(register__n13347), .Y(register__n2288) );
  INVx1_ASAP7_75t_R register___U6148 ( .A(register__n13336), .Y(register__n2289) );
  HB1xp67_ASAP7_75t_R register___U6149 ( .A(register__n12891), .Y(register__n3689) );
  HB1xp67_ASAP7_75t_R register___U6150 ( .A(register__n12890), .Y(register__n3333) );
  HB1xp67_ASAP7_75t_R register___U6151 ( .A(register__n12907), .Y(register__n2988) );
  INVx1_ASAP7_75t_R register___U6152 ( .A(register__n13335), .Y(register__n2290) );
  INVx1_ASAP7_75t_R register___U6153 ( .A(register__n13341), .Y(register__n2291) );
  INVx1_ASAP7_75t_R register___U6154 ( .A(register__n13188), .Y(register__n2292) );
  BUFx6f_ASAP7_75t_R register___U6155 ( .A(register__n11734), .Y(register__n4374) );
  INVx1_ASAP7_75t_R register___U6156 ( .A(register__n13351), .Y(register__n2293) );
  INVx1_ASAP7_75t_R register___U6157 ( .A(register__n13355), .Y(register__n2294) );
  INVx1_ASAP7_75t_R register___U6158 ( .A(register__n13350), .Y(register__n2295) );
  INVx1_ASAP7_75t_R register___U6159 ( .A(register__n13354), .Y(register__n2296) );
  INVx1_ASAP7_75t_R register___U6160 ( .A(register__n12702), .Y(register__n2297) );
  INVx2_ASAP7_75t_R register___U6161 ( .A(register__n6804), .Y(register__n9170) );
  CKINVDCx10_ASAP7_75t_R register___U6162 ( .A(register__n11909), .Y(register__n11829) );
  NOR2x1_ASAP7_75t_R register___U6163 ( .A(register__n2298), .B(register__n2299), .Y(register__net35929) );
  NOR2x1_ASAP7_75t_R register___U6164 ( .A(register__n2300), .B(register__n2301), .Y(register__net35927) );
  NAND2xp5_ASAP7_75t_R register___U6165 ( .A(register__n2302), .B(register__n2303), .Y(register__net119141) );
  INVx2_ASAP7_75t_R register___U6166 ( .A(register__net63278), .Y(register__net63246) );
  NAND2x1p5_ASAP7_75t_R register___U6167 ( .A(register__n2304), .B(register__n118), .Y(register__n2302) );
  NAND2x1p5_ASAP7_75t_R register___U6168 ( .A(register__net63278), .B(register__n1183), .Y(register__n2303) );
  NOR2x1p5_ASAP7_75t_R register___U6169 ( .A(register__n1187), .B(register__net97213), .Y(register__n2300) );
  NOR2x2_ASAP7_75t_R register___U6170 ( .A(register__net63162), .B(register__n120), .Y(register__n2301) );
  NOR2x1p5_ASAP7_75t_R register___U6171 ( .A(register__n1569), .B(register__net62994), .Y(register__n2298) );
  NOR2x1p5_ASAP7_75t_R register___U6172 ( .A(register__net106156), .B(register__n1184), .Y(register__n2299) );
  INVx3_ASAP7_75t_R register___U6173 ( .A(register__net97161), .Y(register__n2304) );
  NOR2x1_ASAP7_75t_R register___U6174 ( .A(register__n2311), .B(register__n1888), .Y(register__net36437) );
  NOR2x1_ASAP7_75t_R register___U6175 ( .A(register__n2313), .B(register__n2314), .Y(register__net36418) );
  NAND2xp5_ASAP7_75t_R register___U6176 ( .A(register__n2315), .B(register__n2316), .Y(register__net111561) );
  INVx1_ASAP7_75t_R register___U6177 ( .A(register__n2317), .Y(register__n2316) );
  NAND2x1p5_ASAP7_75t_R register___U6178 ( .A(register__n2318), .B(register__n117), .Y(register__n2315) );
  NOR2x1p5_ASAP7_75t_R register___U6179 ( .A(register__net97245), .B(register__n1659), .Y(register__n2313) );
  NOR2x1p5_ASAP7_75t_R register___U6180 ( .A(register__n106), .B(register__net64690), .Y(register__n2307) );
  NOR2x1p5_ASAP7_75t_R register___U6181 ( .A(register__n111), .B(register__net63346), .Y(register__n2311) );
  NOR2x1p5_ASAP7_75t_R register___U6182 ( .A(register__n114), .B(register__net63010), .Y(register__n2309) );
  NOR2x1p5_ASAP7_75t_R register___U6183 ( .A(register__n110), .B(register__net62674), .Y(register__n2305) );
  INVx3_ASAP7_75t_R register___U6184 ( .A(register__net91523), .Y(register__n2318) );
  NOR2x1p5_ASAP7_75t_R register___U6185 ( .A(register__n116), .B(register__net64858), .Y(register__n2317) );
  A2O1A1Ixp33_ASAP7_75t_R register___U6186 ( .A1(register__n2319), .A2(register__n2320), .B(register__n54), .C(register__n18), 
        .Y(read_reg_data_1[5]) );
  NOR2x1_ASAP7_75t_R register___U6187 ( .A(register__n2325), .B(register__n1865), .Y(register__n2327) );
  NOR2x1_ASAP7_75t_R register___U6188 ( .A(register__n2336), .B(register__n388), .Y(register__n2337) );
  NOR2x1_ASAP7_75t_R register___U6189 ( .A(register__n2341), .B(register__n2342), .Y(register__n2343) );
  NOR3xp33_ASAP7_75t_R register___U6190 ( .A(register__n2349), .B(register__n2324), .C(register__n2327), .Y(register__n2350) );
  OAI211xp5_ASAP7_75t_R register___U6191 ( .A1(register__C6422_net59703), .A2(register__n1978), .B(register__n2346), 
        .C(register__n2350), .Y(register__n2351) );
  OAI21xp5_ASAP7_75t_R register___U6192 ( .A1(register__n2326), .A2(register__n41), .B(register__n2353), .Y(register__n2352) );
  OAI211xp5_ASAP7_75t_R register___U6193 ( .A1(register__net127380), .A2(register__n2328), .B(register__n2354), .C(
        n2355), .Y(register__n2357) );
  OAI211xp5_ASAP7_75t_R register___U6194 ( .A1(register__n2338), .A2(register__n327), .B(register__n2360), .C(register__n2361), 
        .Y(register__n2363) );
  OAI211xp5_ASAP7_75t_R register___U6195 ( .A1(register__n2344), .A2(register__n169), .B(register__n2366), .C(register__n2364), 
        .Y(register__n2365) );
  INVx4_ASAP7_75t_R register___U6196 ( .A(register__net96610), .Y(register__C6423_net60623) );
  INVx3_ASAP7_75t_R register___U6197 ( .A(register__net90077), .Y(register__n2329) );
  INVx2_ASAP7_75t_R register___U6198 ( .A(register__net89861), .Y(register__n2328) );
  INVx2_ASAP7_75t_R register___U6199 ( .A(register__net90109), .Y(register__n2345) );
  INVx2_ASAP7_75t_R register___U6200 ( .A(register__net90037), .Y(register__n2338) );
  AOI21x1_ASAP7_75t_R register___U6201 ( .A1(register__C6422_net70282), .A2(register__net90789), .B(register__n2359), 
        .Y(register__n2360) );
  NOR2x2_ASAP7_75t_R register___U6202 ( .A(register__C6422_net59704), .B(register__C6422_net69762), .Y(register__n2322)
         );
  OAI21x1_ASAP7_75t_R register___U6203 ( .A1(register__n420), .A2(register__n2321), .B(register__n26), .Y(register__n2349) );
  NOR2x1p5_ASAP7_75t_R register___U6204 ( .A(register__net99656), .B(register__n2333), .Y(register__n2335) );
  OAI21x1_ASAP7_75t_R register___U6205 ( .A1(register__n1455), .A2(register__n2334), .B(register__n69), .Y(register__n2359) );
  INVx2_ASAP7_75t_R register___U6206 ( .A(register__net88889), .Y(register__n2321) );
  INVx2_ASAP7_75t_R register___U6207 ( .A(register__net90865), .Y(register__n2325) );
  INVx2_ASAP7_75t_R register___U6208 ( .A(register__net89953), .Y(register__n2326) );
  INVx2_ASAP7_75t_R register___U6209 ( .A(register__net89773), .Y(register__n2332) );
  INVx3_ASAP7_75t_R register___U6210 ( .A(register__net90829), .Y(register__n2333) );
  INVx2_ASAP7_75t_R register___U6211 ( .A(register__net93737), .Y(register__n2344) );
  INVx2_ASAP7_75t_R register___U6212 ( .A(register__net90145), .Y(register__n2334) );
  INVx3_ASAP7_75t_R register___U6213 ( .A(register__net93837), .Y(register__n2331) );
  INVx2_ASAP7_75t_R register___U6214 ( .A(register__net91069), .Y(register__n2341) );
  INVx4_ASAP7_75t_R register___U6215 ( .A(register__net90729), .Y(register__n2336) );
  INVx2_ASAP7_75t_R register___U6216 ( .A(register__net90901), .Y(register__n2339) );
  NOR2x1_ASAP7_75t_R register___U6217 ( .A(register__n2384), .B(register__n1336), .Y(register__n2385) );
  NOR2x1_ASAP7_75t_R register___U6218 ( .A(register__n2390), .B(register__n2342), .Y(register__n2392) );
  NOR2x1_ASAP7_75t_R register___U6219 ( .A(register__n2391), .B(register__n1509), .Y(register__n2393) );
  OAI211xp5_ASAP7_75t_R register___U6220 ( .A1(register__n420), .A2(register__n2371), .B(register__n25), .C(register__n16), .Y(
        n2396) );
  NAND2xp5_ASAP7_75t_R register___U6221 ( .A(register__n2404), .B(register__n2403), .Y(register__n2405) );
  AOI211xp5_ASAP7_75t_R register___U6222 ( .A1(register__net126316), .A2(register__net91001), .B(register__n2405), .C(
        n2406), .Y(register__n2408) );
  OAI211xp5_ASAP7_75t_R register___U6223 ( .A1(register__n2389), .A2(register__n1420), .B(register__n1893), .C(register__n2408), 
        .Y(register__n2410) );
  INVx4_ASAP7_75t_R register___U6224 ( .A(register__net91495), .Y(register__C6422_net59726) );
  INVx4_ASAP7_75t_R register___U6225 ( .A(register__net91527), .Y(register__C6422_net59730) );
  INVx4_ASAP7_75t_R register___U6226 ( .A(register__net91447), .Y(register__C6422_net59731) );
  INVx2_ASAP7_75t_R register___U6227 ( .A(register__net90113), .Y(register__n2389) );
  INVx2_ASAP7_75t_R register___U6228 ( .A(register__net91073), .Y(register__n2390) );
  AOI21x1_ASAP7_75t_R register___U6229 ( .A1(register__net129746), .A2(register__net90793), .B(register__n2385), .Y(
        n2404) );
  INVx2_ASAP7_75t_R register___U6230 ( .A(register__net90041), .Y(register__n2386) );
  INVx2_ASAP7_75t_R register___U6231 ( .A(register__net89913), .Y(register__n2391) );
  NOR2x1p5_ASAP7_75t_R register___U6232 ( .A(register__n1455), .B(register__n2382), .Y(register__n2383) );
  NOR2x1p5_ASAP7_75t_R register___U6233 ( .A(register__net109643), .B(register__n2378), .Y(register__n2380) );
  INVx2_ASAP7_75t_R register___U6234 ( .A(register__net89817), .Y(register__n2384) );
  INVx3_ASAP7_75t_R register___U6235 ( .A(register__net90149), .Y(register__n2382) );
  INVx2_ASAP7_75t_R register___U6236 ( .A(register__net90905), .Y(register__n2387) );
  INVx2_ASAP7_75t_R register___U6237 ( .A(register__net88893), .Y(register__n2371) );
  INVx2_ASAP7_75t_R register___U6238 ( .A(register__net89865), .Y(register__n2376) );
  INVx3_ASAP7_75t_R register___U6239 ( .A(register__net90081), .Y(register__n2378) );
  INVx2_ASAP7_75t_R register___U6240 ( .A(register__net90833), .Y(register__n2381) );
  NOR2x1p5_ASAP7_75t_R register___U6241 ( .A(register__n66), .B(register__n2370), .Y(register__n2374) );
  INVx3_ASAP7_75t_R register___U6242 ( .A(register__net91463), .Y(register__n2370) );
  INVx2_ASAP7_75t_R register___U6243 ( .A(register__net90937), .Y(register__n2377) );
  NOR2x1_ASAP7_75t_R register___U6244 ( .A(register__n2416), .B(register__n1180), .Y(register__n2417) );
  NOR2x1_ASAP7_75t_R register___U6245 ( .A(register__n2418), .B(register__n2419), .Y(register__n2421) );
  NAND3xp33_ASAP7_75t_R register___U6246 ( .A(register__n2440), .B(register__n2441), .C(register__n2438), .Y(register__n2439) );
  NOR2x1_ASAP7_75t_R register___U6247 ( .A(register__n2421), .B(register__n2422), .Y(register__n2440) );
  NOR4xp75_ASAP7_75t_R register___U6248 ( .A(register__n2426), .B(register__n78), .C(register__n2425), .D(register__n1899), .Y(
        n2448) );
  OAI211xp5_ASAP7_75t_R register___U6249 ( .A1(register__n2436), .A2(register__n_cell_125074_net170554), .B(
        n2455), .C(register__n2456), .Y(register__n2454) );
  AO21x1_ASAP7_75t_R register___U6250 ( .A1(register__n927), .A2(register__net93464), .B(register__n2454), .Y(register__n2457) );
  AO21x1_ASAP7_75t_R register___U6251 ( .A1(register__n642), .A2(register__net90017), .B(register__n2457), .Y(register__n2458) );
  INVx1_ASAP7_75t_R register___U6252 ( .A(register__net107815), .Y(register__n2460) );
  OAI211xp5_ASAP7_75t_R register___U6253 ( .A1(register__n1439), .A2(register__n2414), .B(register__n2459), .C(register__n2442), 
        .Y(register__n2461) );
  INVx1_ASAP7_75t_R register___U6254 ( .A(register__n2429), .Y(register__n2449) );
  NAND2xp5_ASAP7_75t_R register___U6255 ( .A(register__n2462), .B(register__n2461), .Y(register__n2412) );
  INVx4_ASAP7_75t_R register___U6256 ( .A(register__net88977), .Y(register__C6422_net60224) );
  INVx2_ASAP7_75t_R register___U6257 ( .A(register__net88957), .Y(register__C6423_net61141) );
  INVx2_ASAP7_75t_R register___U6258 ( .A(register__net89889), .Y(register__n2414) );
  INVx2_ASAP7_75t_R register___U6259 ( .A(register__net88913), .Y(register__n2423) );
  NOR2x1p5_ASAP7_75t_R register___U6260 ( .A(register__n277), .B(register__n2420), .Y(register__n2422) );
  NOR2x1p5_ASAP7_75t_R register___U6261 ( .A(register__net126725), .B(register__n2413), .Y(register__n2415) );
  INVx2_ASAP7_75t_R register___U6262 ( .A(register__net90853), .Y(register__n2427) );
  INVx2_ASAP7_75t_R register___U6263 ( .A(register__net93853), .Y(register__n2418) );
  INVx6_ASAP7_75t_R register___U6264 ( .A(register__net89793), .Y(register__n2420) );
  INVx2_ASAP7_75t_R register___U6265 ( .A(register__net96903), .Y(register__n2416) );
  INVx3_ASAP7_75t_R register___U6266 ( .A(register__net106940), .Y(register__n2413) );
  INVx2_ASAP7_75t_R register___U6267 ( .A(register__net90813), .Y(register__n2433) );
  INVx4_ASAP7_75t_R register___U6268 ( .A(register__net91021), .Y(register__n2430) );
  INVx4_ASAP7_75t_R register___U6269 ( .A(register__net90761), .Y(register__n2431) );
  INVx2_ASAP7_75t_R register___U6270 ( .A(register__net93420), .Y(register__n2436) );
  NOR2x1p5_ASAP7_75t_R register___U6271 ( .A(register__net130031), .B(register__n2428), .Y(register__n2429) );
  INVx4_ASAP7_75t_R register___U6272 ( .A(register__net89845), .Y(register__n2432) );
  INVx3_ASAP7_75t_R register___U6273 ( .A(register__net90169), .Y(register__n2428) );
  INVx2_ASAP7_75t_R register___U6274 ( .A(register__net93440), .Y(register__n2434) );
  NOR3xp33_ASAP7_75t_R register___U6275 ( .A(register__n2464), .B(register__n2465), .C(register__n2466), .Y(register__n2463) );
  NOR2x1_ASAP7_75t_R register___U6276 ( .A(register__n2474), .B(register__n_cell_124679_net155998), .Y(register__n2476)
         );
  NOR2x1_ASAP7_75t_R register___U6277 ( .A(register__n2478), .B(register__n_cell_124679_net156005), .Y(register__n2480)
         );
  NOR2x1_ASAP7_75t_R register___U6278 ( .A(register__n2481), .B(register__n_cell_124679_net155985), .Y(register__n2482)
         );
  NOR2x1_ASAP7_75t_R register___U6279 ( .A(register__n2487), .B(register__n1179), .Y(register__n2488) );
  NOR2x1_ASAP7_75t_R register___U6280 ( .A(register__n2496), .B(register__n453), .Y(register__n2497) );
  NOR2x1_ASAP7_75t_R register___U6281 ( .A(register__net150875), .B(register__n2498), .Y(register__n2499) );
  NOR3xp33_ASAP7_75t_R register___U6282 ( .A(register__n2501), .B(register__n2471), .C(register__n2472), .Y(register__n2503) );
  NOR2x1_ASAP7_75t_R register___U6283 ( .A(register__n2475), .B(register__n2476), .Y(register__n2504) );
  NOR2x1_ASAP7_75t_R register___U6284 ( .A(register__n2479), .B(register__n2480), .Y(register__n2505) );
  NAND3xp33_ASAP7_75t_R register___U6285 ( .A(register__n2505), .B(register__n2504), .C(register__n2503), .Y(register__n2465) );
  NOR2x1_ASAP7_75t_R register___U6286 ( .A(register__n1891), .B(register__n2495), .Y(register__n2515) );
  NAND3xp33_ASAP7_75t_R register___U6287 ( .A(register__n2520), .B(register__n2521), .C(register__n2522), .Y(register__n2519) );
  OAI211xp5_ASAP7_75t_R register___U6288 ( .A1(register__n2013), .A2(register__n2493), .B(register__n2515), .C(register__n2523), 
        .Y(register__n2466) );
  INVx1_ASAP7_75t_R register___U6289 ( .A(register__n2499), .Y(register__n2521) );
  INVx1_ASAP7_75t_R register___U6290 ( .A(register__n2500), .Y(register__n2467) );
  INVx4_ASAP7_75t_R register___U6291 ( .A(register__net103926), .Y(register__C6422_net59832) );
  INVx4_ASAP7_75t_R register___U6292 ( .A(register__net97177), .Y(register__C6423_net60748) );
  INVx4_ASAP7_75t_R register___U6293 ( .A(register__net91219), .Y(register__C6423_net60749) );
  AOI21x1_ASAP7_75t_R register___U6294 ( .A1(register__net90397), .A2(register__net139572), .B(register__n2482), .Y(
        n2506) );
  INVx2_ASAP7_75t_R register___U6295 ( .A(register__net88821), .Y(register__n2493) );
  NOR2x1p5_ASAP7_75t_R register___U6296 ( .A(register__net122247), .B(register__n2477), .Y(register__n2479) );
  NOR2x1p5_ASAP7_75t_R register___U6297 ( .A(register__net99872), .B(register__n2473), .Y(register__n2475) );
  OAI21x1_ASAP7_75t_R register___U6298 ( .A1(register__net99861), .A2(register__n2468), .B(register__n2502), .Y(register__n2501)
         );
  NOR2x2_ASAP7_75t_R register___U6299 ( .A(register__C6423_net60748), .B(register__net107119), .Y(register__n2495) );
  INVx2_ASAP7_75t_R register___U6300 ( .A(register__net89281), .Y(register__n2481) );
  INVx3_ASAP7_75t_R register___U6301 ( .A(register__net89205), .Y(register__n2490) );
  INVx2_ASAP7_75t_R register___U6302 ( .A(register__net93805), .Y(register__n2489) );
  INVx3_ASAP7_75t_R register___U6303 ( .A(register__net104579), .Y(register__n2483) );
  INVx2_ASAP7_75t_R register___U6304 ( .A(register__net89289), .Y(register__n2484) );
  INVx3_ASAP7_75t_R register___U6305 ( .A(register__net90649), .Y(register__n2477) );
  INVx2_ASAP7_75t_R register___U6306 ( .A(register__net89213), .Y(register__n2478) );
  INVx3_ASAP7_75t_R register___U6307 ( .A(register__net90405), .Y(register__n2473) );
  INVx2_ASAP7_75t_R register___U6308 ( .A(register__net89461), .Y(register__n2474) );
  INVx2_ASAP7_75t_R register___U6309 ( .A(register__net89273), .Y(register__n2468) );
  INVx4_ASAP7_75t_R register___U6310 ( .A(register__net90457), .Y(register__n2469) );
  INVx6_ASAP7_75t_R register___U6311 ( .A(register__net89209), .Y(register__n2470) );
  NAND2x1p5_ASAP7_75t_R register___U6312 ( .A(register__net110413), .B(register__net96863), .Y(register__n2518) );
  NAND2x1p5_ASAP7_75t_R register___U6313 ( .A(register__net137463), .B(register__net88404), .Y(register__n2520) );
  INVx2_ASAP7_75t_R register___U6314 ( .A(register__net90393), .Y(register__n2487) );
  INVx4_ASAP7_75t_R register___U6315 ( .A(register__net89285), .Y(register__n2496) );
  INVx2_ASAP7_75t_R register___U6316 ( .A(register__net93404), .Y(register__n2498) );
  INVx2_ASAP7_75t_R register___U6317 ( .A(register__net105530), .Y(register__n2524) );
  A2O1A1Ixp33_ASAP7_75t_R register___U6318 ( .A1(register__n2527), .A2(register__n2528), .B(register__n1949), .C(register__n2529), 
        .Y(read_reg_data_2[29]) );
  NOR2x1_ASAP7_75t_R register___U6319 ( .A(register__net150043), .B(register__n2536), .Y(register__n2538) );
  NOR2x1_ASAP7_75t_R register___U6320 ( .A(register__n2540), .B(register__n_cell_124938_net165675), .Y(register__n2542)
         );
  NOR2x1_ASAP7_75t_R register___U6321 ( .A(register__n2546), .B(register__n_cell_125074_net170535), .Y(register__n2547)
         );
  NOR2x1_ASAP7_75t_R register___U6322 ( .A(register__n2548), .B(register__n1873), .Y(register__n2549) );
  NOR2x1_ASAP7_75t_R register___U6323 ( .A(register__n2550), .B(register__n276), .Y(register__n2551) );
  NOR2x1_ASAP7_75t_R register___U6324 ( .A(register__n2555), .B(register__n435), .Y(register__n2556) );
  NOR2x1_ASAP7_75t_R register___U6325 ( .A(register__n2564), .B(register__n2538), .Y(register__n2563) );
  OAI21xp5_ASAP7_75t_R register___U6326 ( .A1(register__n2013), .A2(register__n2531), .B(register__n2560), .Y(register__n2565) );
  OAI211xp5_ASAP7_75t_R register___U6327 ( .A1(register__n1903), .A2(register__n2541), .B(register__n2567), .C(register__n2568), 
        .Y(register__n2566) );
  NOR3xp33_ASAP7_75t_R register___U6328 ( .A(register__n2569), .B(register__n2547), .C(register__n2549), .Y(register__n2567) );
  OAI21xp5_ASAP7_75t_R register___U6329 ( .A1(register__n2553), .A2(register__n_cell_125074_net170554), .B(
        n2574), .Y(register__n2573) );
  AOI211xp5_ASAP7_75t_R register___U6330 ( .A1(register__n642), .A2(register__net89013), .B(register__n2577), .C(register__n2571), 
        .Y(register__n2576) );
  OAI211xp5_ASAP7_75t_R register___U6331 ( .A1(register__n277), .A2(register__n2557), .B(register__n2579), .C(register__n2580), 
        .Y(register__n2577) );
  OAI211xp5_ASAP7_75t_R register___U6332 ( .A1(register__C6423_net72242), .A2(register__n2554), .B(register__n2575), 
        .C(register__n2576), .Y(register__n2581) );
  INVx1_ASAP7_75t_R register___U6333 ( .A(register__n2582), .Y(register__n2561) );
  INVx1_ASAP7_75t_R register___U6334 ( .A(register__n2583), .Y(register__n2564) );
  INVx1_ASAP7_75t_R register___U6335 ( .A(register__n2558), .Y(register__n2529) );
  INVx4_ASAP7_75t_R register___U6336 ( .A(register__net91203), .Y(register__C6423_net61245) );
  NAND2x1p5_ASAP7_75t_R register___U6337 ( .A(register__net91045), .B(register__C6423_net61318), .Y(register__n2584) );
  INVx2_ASAP7_75t_R register___U6338 ( .A(register__net90233), .Y(register__n2554) );
  INVx2_ASAP7_75t_R register___U6339 ( .A(register__net89445), .Y(register__n2541) );
  INVx4_ASAP7_75t_R register___U6340 ( .A(register__net88764), .Y(register__n2531) );
  OAI21x1_ASAP7_75t_R register___U6341 ( .A1(register__net122250), .A2(register__n2545), .B(register__n76), .Y(register__n2569)
         );
  INVx2_ASAP7_75t_R register___U6342 ( .A(register__net89441), .Y(register__n2553) );
  NAND2x1p5_ASAP7_75t_R register___U6343 ( .A(register__net89001), .B(register__n1906), .Y(register__n2574) );
  INVx2_ASAP7_75t_R register___U6344 ( .A(register__net93408), .Y(register__n2557) );
  INVx2_ASAP7_75t_R register___U6345 ( .A(register__net93673), .Y(register__n2552) );
  INVx2_ASAP7_75t_R register___U6346 ( .A(register__net96843), .Y(register__n2545) );
  INVx2_ASAP7_75t_R register___U6347 ( .A(register__net91583), .Y(register__n2546) );
  INVx2_ASAP7_75t_R register___U6348 ( .A(register__net96915), .Y(register__n2548) );
  INVx4_ASAP7_75t_R register___U6349 ( .A(register__net88756), .Y(register__n2532) );
  INVx3_ASAP7_75t_R register___U6350 ( .A(register__net90629), .Y(register__n2543) );
  INVx3_ASAP7_75t_R register___U6351 ( .A(register__net88997), .Y(register__n2537) );
  INVx2_ASAP7_75t_R register___U6352 ( .A(register__net90221), .Y(register__n2540) );
  INVx6_ASAP7_75t_R register___U6353 ( .A(register__net88760), .Y(register__n2530) );
  INVx2_ASAP7_75t_R register___U6354 ( .A(register__net89005), .Y(register__n2555) );
  INVx2_ASAP7_75t_R register___U6355 ( .A(register__net90213), .Y(register__n2550) );
  INVx2_ASAP7_75t_R register___U6356 ( .A(register__net90237), .Y(register__n2536) );
  NOR3xp33_ASAP7_75t_R register___U6357 ( .A(register__n2586), .B(register__n2587), .C(register__n2588), .Y(register__n2585) );
  NOR2x1_ASAP7_75t_R register___U6358 ( .A(register__n2596), .B(register__n1181), .Y(register__n2597) );
  NOR2x1_ASAP7_75t_R register___U6359 ( .A(register__net150043), .B(register__n2599), .Y(register__n2601) );
  NOR2x1_ASAP7_75t_R register___U6360 ( .A(register__n2602), .B(register__n_cell_124938_net165675), .Y(register__n2604)
         );
  NOR2x1_ASAP7_75t_R register___U6361 ( .A(register__n2607), .B(register__n_cell_125074_net170535), .Y(register__n2608)
         );
  NOR2x1_ASAP7_75t_R register___U6362 ( .A(register__n2609), .B(register__n276), .Y(register__n2610) );
  NOR2x1_ASAP7_75t_R register___U6363 ( .A(register__n2597), .B(register__n2595), .Y(register__n2621) );
  OAI211xp5_ASAP7_75t_R register___U6364 ( .A1(register__n2013), .A2(register__n2590), .B(register__n2620), .C(register__n2623), 
        .Y(register__n2586) );
  AO21x1_ASAP7_75t_R register___U6365 ( .A1(register__net137463), .A2(register__net90661), .B(register__n2608), .Y(
        n2626) );
  OAI211xp5_ASAP7_75t_R register___U6366 ( .A1(register__net130030), .A2(register__n2600), .B(register__n2624), .C(
        n2628), .Y(register__n2587) );
  AO21x1_ASAP7_75t_R register___U6367 ( .A1(register__n2022), .A2(register__net89613), .B(register__n2610), .Y(register__n2629)
         );
  AOI21xp5_ASAP7_75t_R register___U6368 ( .A1(register__C6423_net74857), .A2(register__net89589), .B(register__n2629), 
        .Y(register__n2630) );
  OAI211xp5_ASAP7_75t_R register___U6369 ( .A1(register__n2613), .A2(register__n1650), .B(register__n2632), .C(register__n2630), 
        .Y(register__n2631) );
  INVx1_ASAP7_75t_R register___U6370 ( .A(register__n2614), .Y(register__n2589) );
  INVx2_ASAP7_75t_R register___U6371 ( .A(register__net91375), .Y(register__C6422_net59856) );
  INVx2_ASAP7_75t_R register___U6372 ( .A(register__net106200), .Y(register__C6422_net59860) );
  INVx4_ASAP7_75t_R register___U6373 ( .A(register__net91347), .Y(register__C6423_net60775) );
  INVx4_ASAP7_75t_R register___U6374 ( .A(register__net91367), .Y(register__C6423_net60777) );
  INVx2_ASAP7_75t_R register___U6375 ( .A(register__net88885), .Y(register__n2590) );
  INVx2_ASAP7_75t_R register___U6376 ( .A(register__net89593), .Y(register__n2600) );
  INVx4_ASAP7_75t_R register___U6377 ( .A(register__net90673), .Y(register__n2605) );
  INVx2_ASAP7_75t_R register___U6378 ( .A(register__net89673), .Y(register__n2603) );
  OAI21x1_ASAP7_75t_R register___U6379 ( .A1(register__net122250), .A2(register__n2606), .B(register__n2627), .Y(register__n2625)
         );
  INVx6_ASAP7_75t_R register___U6380 ( .A(register__net88512), .Y(register__n2594) );
  INVx2_ASAP7_75t_R register___U6381 ( .A(register__net89617), .Y(register__n2592) );
  INVx2_ASAP7_75t_R register___U6382 ( .A(register__net93817), .Y(register__n2598) );
  INVx2_ASAP7_75t_R register___U6383 ( .A(register__net90677), .Y(register__n2602) );
  INVx4_ASAP7_75t_R register___U6384 ( .A(register__net90713), .Y(register__n2606) );
  INVx2_ASAP7_75t_R register___U6385 ( .A(register__net90681), .Y(register__n2613) );
  INVx2_ASAP7_75t_R register___U6386 ( .A(register__net105518), .Y(register__n2633) );
  INVx4_ASAP7_75t_R register___U6387 ( .A(register__net89657), .Y(register__n2607) );
  INVx2_ASAP7_75t_R register___U6388 ( .A(register__net90657), .Y(register__n2596) );
  INVx3_ASAP7_75t_R register___U6389 ( .A(register__net88604), .Y(register__n2593) );
  INVx4_ASAP7_75t_R register___U6390 ( .A(register__net90669), .Y(register__n2599) );
  INVx4_ASAP7_75t_R register___U6391 ( .A(register__net89597), .Y(register__n2611) );
  INVx4_ASAP7_75t_R register___U6392 ( .A(register__net90717), .Y(register__n2609) );
  NOR2x1_ASAP7_75t_R register___U6393 ( .A(register__n2645), .B(register__n260), .Y(register__n2647) );
  NOR2x1_ASAP7_75t_R register___U6394 ( .A(register__n2652), .B(register__n327), .Y(register__n2653) );
  OAI21xp5_ASAP7_75t_R register___U6395 ( .A1(register__n2641), .A2(register__n1864), .B(register__n2663), .Y(register__n2662) );
  NOR2x1_ASAP7_75t_R register___U6396 ( .A(register__n2640), .B(register__n2639), .Y(register__n2663) );
  NOR3xp33_ASAP7_75t_R register___U6397 ( .A(register__n2660), .B(register__n2662), .C(register__n2661), .Y(register__n2664) );
  OAI21xp5_ASAP7_75t_R register___U6398 ( .A1(register__n2643), .A2(register__n_cell_124812_net160756), .B(
        n2667), .Y(register__n2666) );
  OAI211xp5_ASAP7_75t_R register___U6399 ( .A1(register__net127380), .A2(register__n2642), .B(register__n2668), .C(
        n2671), .Y(register__n2672) );
  OAI211xp5_ASAP7_75t_R register___U6400 ( .A1(register__n2654), .A2(register__n2342), .B(register__n2678), .C(register__n2675), 
        .Y(register__n2677) );
  OAI211xp5_ASAP7_75t_R register___U6401 ( .A1(register__n2651), .A2(register__C6422_net59572), .B(register__n2673), 
        .C(register__n2676), .Y(register__n2685) );
  INVx4_ASAP7_75t_R register___U6402 ( .A(register__net91263), .Y(register__C6423_net61114) );
  INVx2_ASAP7_75t_R register___U6403 ( .A(register__net90637), .Y(register__n2651) );
  INVx2_ASAP7_75t_R register___U6404 ( .A(register__net90265), .Y(register__n2658) );
  INVx2_ASAP7_75t_R register___U6405 ( .A(register__net90249), .Y(register__n2654) );
  INVx2_ASAP7_75t_R register___U6406 ( .A(register__net89649), .Y(register__n2652) );
  INVx2_ASAP7_75t_R register___U6407 ( .A(register__net88861), .Y(register__n2638) );
  INVx2_ASAP7_75t_R register___U6408 ( .A(register__net89053), .Y(register__n2642) );
  OAI21x1_ASAP7_75t_R register___U6409 ( .A1(register__net109844), .A2(register__n2636), .B(register__n23), .Y(register__n2660)
         );
  INVx2_ASAP7_75t_R register___U6410 ( .A(register__net88504), .Y(register__n2656) );
  AOI21x1_ASAP7_75t_R register___U6411 ( .A1(register__C6422_net70534), .A2(register__net89049), .B(register__n2657), 
        .Y(register__n2679) );
  INVx4_ASAP7_75t_R register___U6412 ( .A(register__net90257), .Y(register__n2650) );
  INVx2_ASAP7_75t_R register___U6413 ( .A(register__net89037), .Y(register__n2649) );
  INVx4_ASAP7_75t_R register___U6414 ( .A(register__net88785), .Y(register__n2636) );
  INVx2_ASAP7_75t_R register___U6415 ( .A(register__net90541), .Y(register__n2641) );
  INVx4_ASAP7_75t_R register___U6416 ( .A(register__net90537), .Y(register__n2643) );
  INVx2_ASAP7_75t_R register___U6417 ( .A(register__net90545), .Y(register__n2648) );
  NOR2x2_ASAP7_75t_R register___U6418 ( .A(register__net105510), .B(register__n802), .Y(register__n2640) );
  NOR2x1p5_ASAP7_75t_R register___U6419 ( .A(register__n1398), .B(register__n2644), .Y(register__n2646) );
  INVx4_ASAP7_75t_R register___U6420 ( .A(register__net88416), .Y(register__n2655) );
  INVx6_ASAP7_75t_R register___U6421 ( .A(register__net91331), .Y(register__n2635) );
  INVx3_ASAP7_75t_R register___U6422 ( .A(register__net91335), .Y(register__n2637) );
  INVx2_ASAP7_75t_R register___U6423 ( .A(register__net89417), .Y(register__n2645) );
  INVx3_ASAP7_75t_R register___U6424 ( .A(register__net93793), .Y(register__n2644) );
  NOR2x1_ASAP7_75t_R register___U6425 ( .A(register__n2712), .B(register__n454), .Y(register__n2714) );
  NOR2x1_ASAP7_75t_R register___U6426 ( .A(register__n2019), .B(register__n2715), .Y(register__n2716) );
  OAI221xp5_ASAP7_75t_R register___U6427 ( .A1(register__net94610), .A2(register__net107119), .B1(
        C6422_net59961), .B2(register__n710), .C(register__n2721), .Y(register__n2722) );
  AO21x1_ASAP7_75t_R register___U6428 ( .A1(register__net125170), .A2(register__net88412), .B(register__n2697), .Y(
        n2723) );
  NOR2x1_ASAP7_75t_R register___U6429 ( .A(register__n2723), .B(register__n2694), .Y(register__n2724) );
  OAI21xp5_ASAP7_75t_R register___U6430 ( .A1(register__C6423_net72245), .A2(register__n2698), .B(register__n2726), .Y(
        n2728) );
  OAI211xp5_ASAP7_75t_R register___U6431 ( .A1(register__n112), .A2(register__n2704), .B(register__n2731), .C(register__n2732), 
        .Y(register__n2730) );
  AO21x1_ASAP7_75t_R register___U6432 ( .A1(register__net137463), .A2(register__net90521), .B(register__n2714), .Y(
        n2734) );
  AO21x1_ASAP7_75t_R register___U6433 ( .A1(register__n924), .A2(register__net93713), .B(register__n2734), .Y(register__n2735) );
  OAI21xp5_ASAP7_75t_R register___U6434 ( .A1(register__n2717), .A2(register__n2437), .B(register__n2736), .Y(register__n2737) );
  NAND2xp5_ASAP7_75t_R register___U6435 ( .A(register__n2729), .B(register__n2738), .Y(register__n2688) );
  INVx1_ASAP7_75t_R register___U6436 ( .A(register__n2718), .Y(register__n2689) );
  INVx2_ASAP7_75t_R register___U6437 ( .A(register__net93576), .Y(register__C6422_net59965) );
  INVx4_ASAP7_75t_R register___U6438 ( .A(register__net103940), .Y(register__C6423_net60880) );
  INVx4_ASAP7_75t_R register___U6439 ( .A(register__net99037), .Y(register__net94610) );
  OAI21x1_ASAP7_75t_R register___U6440 ( .A1(register__n1439), .A2(register__n2696), .B(register__n2724), .Y(register__n2725) );
  INVx2_ASAP7_75t_R register___U6441 ( .A(register__net88584), .Y(register__n2704) );
  NAND2x1p5_ASAP7_75t_R register___U6442 ( .A(register__net102304), .B(register__net90689), .Y(register__n2731) );
  INVx3_ASAP7_75t_R register___U6443 ( .A(register__net89393), .Y(register__n2701) );
  INVx2_ASAP7_75t_R register___U6444 ( .A(register__net91591), .Y(register__n2717) );
  INVx3_ASAP7_75t_R register___U6445 ( .A(register__net91259), .Y(register__n2690) );
  INVx2_ASAP7_75t_R register___U6446 ( .A(register__net89409), .Y(register__n2696) );
  INVx2_ASAP7_75t_R register___U6447 ( .A(register__net90525), .Y(register__n2698) );
  NOR2x1p5_ASAP7_75t_R register___U6448 ( .A(register__n277), .B(register__n2693), .Y(register__n2694) );
  INVx3_ASAP7_75t_R register___U6449 ( .A(register__net90533), .Y(register__n2707) );
  INVx2_ASAP7_75t_R register___U6450 ( .A(register__net88500), .Y(register__n2705) );
  INVx2_ASAP7_75t_R register___U6451 ( .A(register__C6423_net69178), .Y(register__n_cell_124679_net155998) );
  INVx2_ASAP7_75t_R register___U6452 ( .A(register__net89553), .Y(register__n2708) );
  INVx4_ASAP7_75t_R register___U6453 ( .A(register__net90529), .Y(register__n2711) );
  INVx4_ASAP7_75t_R register___U6454 ( .A(register__net89405), .Y(register__n2712) );
  INVx2_ASAP7_75t_R register___U6455 ( .A(register__net89641), .Y(register__n2715) );
  INVx3_ASAP7_75t_R register___U6456 ( .A(register__net96819), .Y(register__n2693) );
  INVx2_ASAP7_75t_R register___U6457 ( .A(register__net93797), .Y(register__n2700) );
  INVx2_ASAP7_75t_R register___U6458 ( .A(register__net89401), .Y(register__n2699) );
  INVx3_ASAP7_75t_R register___U6459 ( .A(register__net104592), .Y(register__n2695) );
  AO22x1_ASAP7_75t_R register___U6460 ( .A1(register__n9871), .A2(register__n481), .B1(register__n10285), .B2(register__n640), 
        .Y(register__n11637) );
  AND3x1_ASAP7_75t_R register___U6461 ( .A(register__n11079), .B(register__n11080), .C(register__n11078), .Y(register__n2768) );
  INVx2_ASAP7_75t_R register___U6462 ( .A(register__n5119), .Y(register__n7672) );
  HB1xp67_ASAP7_75t_R register___U6463 ( .A(register__n11657), .Y(register__n3210) );
  INVxp67_ASAP7_75t_R register___U6464 ( .A(register__n6021), .Y(register__n9206) );
  HB1xp67_ASAP7_75t_R register___U6465 ( .A(register__n6022), .Y(register__n6021) );
  AO22x1_ASAP7_75t_R register___U6466 ( .A1(register__n9780), .A2(register__n85), .B1(register__n10096), .B2(register__n422), .Y(
        n11314) );
  INVxp67_ASAP7_75t_R register___U6467 ( .A(register__net124564), .Y(register__net109574) );
  HB1xp67_ASAP7_75t_R register___U6468 ( .A(register__C6423_net60964), .Y(register__net122897) );
  AO22x1_ASAP7_75t_R register___U6469 ( .A1(register__n9748), .A2(register__n85), .B1(register__n10108), .B2(
        C6423_net61335), .Y(register__n11400) );
  AO22x1_ASAP7_75t_R register___U6470 ( .A1(register__n9802), .A2(register__n85), .B1(register__n10140), .B2(register__n422), .Y(
        n11422) );
  AO22x1_ASAP7_75t_R register___U6471 ( .A1(register__n9897), .A2(register__n85), .B1(register__n10223), .B2(register__n2086), 
        .Y(register__n11672) );
  AO22x1_ASAP7_75t_R register___U6472 ( .A1(register__n9714), .A2(register__net129017), .B1(register__n10044), .B2(
        n2086), .Y(register__n11254) );
  AO22x1_ASAP7_75t_R register___U6473 ( .A1(register__n9774), .A2(register__n85), .B1(register__n10275), .B2(
        C6423_net61335), .Y(register__n11360) );
  INVx2_ASAP7_75t_R register___U6474 ( .A(register__n5108), .Y(register__n7005) );
  INVx2_ASAP7_75t_R register___U6475 ( .A(register__net122896), .Y(register__net100454) );
  AO22x1_ASAP7_75t_R register___U6476 ( .A1(register__n9716), .A2(register__net102299), .B1(register__n10046), .B2(register__n422), .Y(register__n11234) );
  INVx2_ASAP7_75t_R register___U6477 ( .A(register__n12034), .Y(register__n12018) );
  INVx1_ASAP7_75t_R register___U6478 ( .A(register__n11558), .Y(register__n2743) );
  INVxp33_ASAP7_75t_R register___U6479 ( .A(register__n239), .Y(register__net150880) );
  INVxp33_ASAP7_75t_R register___U6480 ( .A(register__net150878), .Y(register__net150882) );
  INVxp33_ASAP7_75t_R register___U6481 ( .A(register__net150878), .Y(register__net150887) );
  HB1xp67_ASAP7_75t_R register___U6482 ( .A(register__n1998), .Y(register__net121558) );
  HB1xp67_ASAP7_75t_R register___U6483 ( .A(register__net124565), .Y(register__net124564) );
  AO22x1_ASAP7_75t_R register___U6484 ( .A1(register__net90681), .A2(register__n38), .B1(register__net89581), .B2(
        C6422_net70678), .Y(register__n10729) );
  HB1xp67_ASAP7_75t_R register___U6485 ( .A(register__n11370), .Y(register__n6022) );
  INVxp67_ASAP7_75t_R register___U6486 ( .A(register__net139811), .Y(register__net122188) );
  HB1xp67_ASAP7_75t_R register___U6487 ( .A(register__net139812), .Y(register__net139811) );
  BUFx12f_ASAP7_75t_R register___U6488 ( .A(register__net67414), .Y(register__net67412) );
  INVx1_ASAP7_75t_R register___U6489 ( .A(register__n12272), .Y(register__n12259) );
  BUFx2_ASAP7_75t_R register___U6490 ( .A(register__n12078), .Y(register__n12070) );
  INVx2_ASAP7_75t_R register___U6491 ( .A(register__n12070), .Y(register__n12057) );
  INVxp33_ASAP7_75t_R register___U6492 ( .A(register__n5264), .Y(register__n5665) );
  INVx6_ASAP7_75t_R register___U6493 ( .A(register__n5074), .Y(register__n8564) );
  HB1xp67_ASAP7_75t_R register___U6494 ( .A(register__n3210), .Y(register__n6719) );
  INVxp67_ASAP7_75t_R register___U6495 ( .A(register__n5258), .Y(register__n8569) );
  AO22x1_ASAP7_75t_R register___U6496 ( .A1(register__n9642), .A2(register__n1909), .B1(register__n9969), .B2(register__n381), 
        .Y(register__n10972) );
  CKINVDCx10_ASAP7_75t_R register___U6497 ( .A(register__n12075), .Y(register__n5074) );
  INVxp33_ASAP7_75t_R register___U6498 ( .A(register__n5556), .Y(register__n7604) );
  HB1xp67_ASAP7_75t_R register___U6499 ( .A(register__n4578), .Y(register__n12272) );
  AND3x1_ASAP7_75t_R register___U6500 ( .A(register__n10657), .B(register__n763), .C(register__n10656), .Y(register__n2776) );
  HB1xp67_ASAP7_75t_R register___U6501 ( .A(register__n11656), .Y(register__n3110) );
  INVxp33_ASAP7_75t_R register___U6502 ( .A(register__n4442), .Y(register__n8267) );
  AO22x1_ASAP7_75t_R register___U6503 ( .A1(register__n8807), .A2(register__n156), .B1(register__n8817), .B2(register__n381), .Y(
        n10949) );
  HB1xp67_ASAP7_75t_R register___U6504 ( .A(register__n10754), .Y(register__n5264) );
  HB1xp67_ASAP7_75t_R register___U6505 ( .A(register__n4443), .Y(register__n4442) );
  AND3x1_ASAP7_75t_R register___U6506 ( .A(register__n11034), .B(register__n11036), .C(register__n11035), .Y(register__n2767) );
  HB1xp67_ASAP7_75t_R register___U6507 ( .A(register__n11637), .Y(register__n3239) );
  AO22x1_ASAP7_75t_R register___U6508 ( .A1(register__net88404), .A2(register__n3), .B1(register__net88496), .B2(register__n281), 
        .Y(register__n10715) );
  AO22x1_ASAP7_75t_R register___U6509 ( .A1(register__n6915), .A2(register__n230), .B1(register__net150889), .B2(register__n9382), 
        .Y(register__n11558) );
  INVx6_ASAP7_75t_R register___U6510 ( .A(register__n12068), .Y(register__n12055) );
  HB1xp67_ASAP7_75t_R register___U6511 ( .A(register__n5259), .Y(register__n5258) );
  AO22x1_ASAP7_75t_R register___U6512 ( .A1(register__n9730), .A2(register__n3), .B1(register__n10098), .B2(register__n233), .Y(
        n10696) );
  AO22x1_ASAP7_75t_R register___U6513 ( .A1(register__n10442), .A2(register__n481), .B1(register__n10426), .B2(
        C6423_net61348), .Y(register__n11656) );
  AO22x1_ASAP7_75t_R register___U6514 ( .A1(register__n9644), .A2(register__n1909), .B1(register__n9971), .B2(register__n381), 
        .Y(register__n10928) );
  HB1xp67_ASAP7_75t_R register___U6515 ( .A(register__n10715), .Y(register__n5556) );
  HB1xp67_ASAP7_75t_R register___U6516 ( .A(register__net36418), .Y(register__net124565) );
  AO22x1_ASAP7_75t_R register___U6517 ( .A1(register__n9879), .A2(register__n1909), .B1(register__n10157), .B2(register__n381), 
        .Y(register__n10754) );
  HB1xp67_ASAP7_75t_R register___U6518 ( .A(register__n10837), .Y(register__n4443) );
  AO22x1_ASAP7_75t_R register___U6519 ( .A1(register__n9658), .A2(register__n156), .B1(register__n9985), .B2(register__n1579), 
        .Y(register__n10546) );
  AO22x1_ASAP7_75t_R register___U6520 ( .A1(register__n9656), .A2(register__n3), .B1(register__n9983), .B2(register__register__n381), .Y(
        n10567) );
  INVxp33_ASAP7_75t_R register___U6521 ( .A(register__n2026), .Y(register__net150060) );
  AND2x2_ASAP7_75t_R register___U6522 ( .A(register__n11720), .B(register__n597), .Y(register__C6423_net61333) );
  HB1xp67_ASAP7_75t_R register___U6523 ( .A(register__C6423_net61333), .Y(register__net98137) );
  AO22x1_ASAP7_75t_R register___U6524 ( .A1(register__net90865), .A2(register__net138040), .B1(register__net89953), 
        .B2(register__C6423_net68766), .Y(register__n11269) );
  AO22x1_ASAP7_75t_R register___U6525 ( .A1(register__n10501), .A2(register__n229), .B1(register__n9246), .B2(register__n1998), 
        .Y(register__n11723) );
  AO22x1_ASAP7_75t_R register___U6526 ( .A1(register__n9676), .A2(register__C6423_net61333), .B1(register__n9419), .B2(
        n767), .Y(register__n11235) );
  BUFx3_ASAP7_75t_R register___U6527 ( .A(register__n11535), .Y(register__n4313) );
  AO22x1_ASAP7_75t_R register___U6528 ( .A1(register__register__n9284), .A2(register__n928), .B1(register__net150892), .B2(register__n10231), .Y(register__n11383) );
  AO22x1_ASAP7_75t_R register___U6529 ( .A1(register__n6924), .A2(register__n883), .B1(register__n6376), .B2(register__net122862), 
        .Y(register__n11713) );
  AO22x1_ASAP7_75t_R register___U6530 ( .A1(register__n12273), .A2(register__n5524), .B1(register__n11845), .B2(register__n11915), 
        .Y(register__n9388) );
  AO22x1_ASAP7_75t_R register___U6531 ( .A1(register__n10493), .A2(register__n883), .B1(register__n7994), .B2(register__net139882), .Y(register__n11332) );
  AO22x1_ASAP7_75t_R register___U6532 ( .A1(register__n9680), .A2(register__net150061), .B1(register__n9927), .B2(register__n767), 
        .Y(register__n11169) );
  AO22x1_ASAP7_75t_R register___U6533 ( .A1(register__n9339), .A2(register__net150059), .B1(register__n9325), .B2(register__n767), 
        .Y(register__n11191) );
  HB1xp67_ASAP7_75t_R register___U6534 ( .A(register__n6033), .Y(register__n5116) );
  AO22x1_ASAP7_75t_R register___U6535 ( .A1(register__n9353), .A2(register__net122579), .B1(register__n8793), .B2(register__n1998), .Y(register__n11654) );
  AO22x1_ASAP7_75t_R register___U6536 ( .A1(register__n9674), .A2(register__n2004), .B1(register__n9921), .B2(register__n2025), 
        .Y(register__n11489) );
  HB1xp67_ASAP7_75t_R register___U6537 ( .A(register__n11397), .Y(register__n5587) );
  BUFx4f_ASAP7_75t_R register___U6538 ( .A(register__n4948), .Y(register__n4947) );
  BUFx3_ASAP7_75t_R register___U6539 ( .A(register__n11058), .Y(register__n4948) );
  BUFx3_ASAP7_75t_R register___U6540 ( .A(register__n11102), .Y(register__n7699) );
  INVx2_ASAP7_75t_R register___U6541 ( .A(register__n5145), .Y(register__n7977) );
  HB1xp67_ASAP7_75t_R register___U6542 ( .A(register__n10696), .Y(register__n5259) );
  AO22x1_ASAP7_75t_R register___U6543 ( .A1(register__n9274), .A2(register__net150048), .B1(register__n10263), .B2(register__n767), .Y(register__n11595) );
  BUFx12f_ASAP7_75t_R register___U6544 ( .A(register__n8562), .Y(register__n3439) );
  INVx2_ASAP7_75t_R register___U6545 ( .A(register__n4947), .Y(register__n8700) );
  BUFx6f_ASAP7_75t_R register___U6546 ( .A(register__net122602), .Y(register__C6423_net72238) );
  AO22x1_ASAP7_75t_R register___U6547 ( .A1(register__n9411), .A2(register__net137440), .B1(register__n9997), .B2(
        C6423_net68764), .Y(register__n11165) );
  BUFx12f_ASAP7_75t_R register___U6548 ( .A(register__n3710), .Y(register__n11873) );
  HB1xp67_ASAP7_75t_R register___U6549 ( .A(register__net94613), .Y(register__net113157) );
  HB1xp67_ASAP7_75t_R register___U6550 ( .A(register__n11587), .Y(register__n5245) );
  NOR2xp33_ASAP7_75t_R register___U6551 ( .A(register__net63998), .B(register__n983), .Y(register__n2750) );
  NOR2xp33_ASAP7_75t_R register___U6552 ( .A(register__net95072), .B(register__n969), .Y(register__n2751) );
  NOR2xp33_ASAP7_75t_R register___U6553 ( .A(register__n2750), .B(register__n2751), .Y(register__n13193) );
  HB1xp67_ASAP7_75t_R register___U6554 ( .A(register__net91591), .Y(register__net95072) );
  HB1xp67_ASAP7_75t_R register___U6555 ( .A(register__n13193), .Y(register__n5782) );
  NOR3xp33_ASAP7_75t_R register___U6556 ( .A(register__n2752), .B(register__n2753), .C(register__n2754), .Y(register__n11521) );
  HB1xp67_ASAP7_75t_R register___U6557 ( .A(register__n11527), .Y(register__n6468) );
  AND3x1_ASAP7_75t_R register___U6558 ( .A(register__n10757), .B(register__n10756), .C(register__n171), .Y(register__n2756) );
  AND2x2_ASAP7_75t_R register___U6559 ( .A(register__n10755), .B(register__n2756), .Y(register__n3720) );
  NOR2xp33_ASAP7_75t_R register___U6560 ( .A(register__n12113), .B(register__n992), .Y(register__n2757) );
  NOR2xp33_ASAP7_75t_R register___U6561 ( .A(register__n10144), .B(register__n973), .Y(register__n2758) );
  NOR2xp33_ASAP7_75t_R register___U6562 ( .A(register__n2757), .B(register__n2758), .Y(register__n13196) );
  HB1xp67_ASAP7_75t_R register___U6563 ( .A(register__n13196), .Y(register__n5778) );
  NOR2xp33_ASAP7_75t_R register___U6564 ( .A(register__n10126), .B(register__n973), .Y(register__n2760) );
  NOR2xp33_ASAP7_75t_R register___U6565 ( .A(register__n99), .B(register__n980), .Y(register__n2761) );
  NOR2xp33_ASAP7_75t_R register___U6566 ( .A(register__n10321), .B(register__n971), .Y(register__n2762) );
  NOR2xp33_ASAP7_75t_R register___U6567 ( .A(register__n2761), .B(register__n2762), .Y(register__n13191) );
  HB1xp67_ASAP7_75t_R register___U6568 ( .A(register__n13191), .Y(register__n5980) );
  NOR2xp33_ASAP7_75t_R register___U6569 ( .A(register__n12282), .B(register__n976), .Y(register__n2763) );
  NOR2xp33_ASAP7_75t_R register___U6570 ( .A(register__n10239), .B(register__n972), .Y(register__n2764) );
  NOR2xp33_ASAP7_75t_R register___U6571 ( .A(register__n2763), .B(register__n2764), .Y(register__n13189) );
  HB1xp67_ASAP7_75t_R register___U6572 ( .A(register__n13189), .Y(register__n5978) );
  AND2x2_ASAP7_75t_R register___U6573 ( .A(register__n7267), .B(register__n11494), .Y(register__n2765) );
  HB1xp67_ASAP7_75t_R register___U6574 ( .A(register__n11495), .Y(register__n7267) );
  AND2x2_ASAP7_75t_R register___U6575 ( .A(register__n8295), .B(register__n2768), .Y(register__n7889) );
  NOR2xp33_ASAP7_75t_R register___U6576 ( .A(register__n10197), .B(register__n975), .Y(register__n2771) );
  HB1xp67_ASAP7_75t_R register___U6577 ( .A(register__n13194), .Y(register__n5975) );
  NOR2xp33_ASAP7_75t_R register___U6578 ( .A(register__n12262), .B(register__n981), .Y(register__n2772) );
  NOR2xp33_ASAP7_75t_R register___U6579 ( .A(register__n10088), .B(register__n970), .Y(register__n2773) );
  NOR2xp33_ASAP7_75t_R register___U6580 ( .A(register__n2772), .B(register__n2773), .Y(register__n13190) );
  HB1xp67_ASAP7_75t_R register___U6581 ( .A(register__n13190), .Y(register__n4402) );
  NOR2xp33_ASAP7_75t_R register___U6582 ( .A(register__n12195), .B(register__n989), .Y(register__n2774) );
  NOR2xp33_ASAP7_75t_R register___U6583 ( .A(register__n10465), .B(register__n974), .Y(register__n2775) );
  NOR2xp33_ASAP7_75t_R register___U6584 ( .A(register__n2774), .B(register__n2775), .Y(register__n13192) );
  HB1xp67_ASAP7_75t_R register___U6585 ( .A(register__n13192), .Y(register__n4067) );
  AND2x2_ASAP7_75t_R register___U6586 ( .A(register__n10655), .B(register__n2776), .Y(register__n8273) );
  AND2x2_ASAP7_75t_R register___U6587 ( .A(register__n5557), .B(register__n2777), .Y(register__n10697) );
  HB1xp67_ASAP7_75t_R register___U6588 ( .A(register__n7604), .Y(register__n5557) );
  AND2x2_ASAP7_75t_R register___U6589 ( .A(register__n5265), .B(register__n2778), .Y(register__n10732) );
  HB1xp67_ASAP7_75t_R register___U6590 ( .A(register__n5665), .Y(register__n5265) );
  HB1xp67_ASAP7_75t_R register___U6591 ( .A(register__n8267), .Y(register__n4444) );
  NOR2xp33_ASAP7_75t_R register___U6592 ( .A(register__n9627), .B(register__n342), .Y(register__n2781) );
  AND2x2_ASAP7_75t_R register___U6593 ( .A(register__n11639), .B(register__n11638), .Y(register__n2784) );
  AND2x2_ASAP7_75t_R register___U6594 ( .A(register__n11679), .B(register__n11678), .Y(register__n2785) );
  AND3x1_ASAP7_75t_R register___U6595 ( .A(register__n2785), .B(register__n11680), .C(register__n2195), .Y(register__n4179) );
  NOR2xp33_ASAP7_75t_R register___U6596 ( .A(register__n10483), .B(register__n215), .Y(register__n2787) );
  AND2x2_ASAP7_75t_R register___U6597 ( .A(register__n9153), .B(register__n2790), .Y(register__n10755) );
  NOR2xp33_ASAP7_75t_R register___U6598 ( .A(register__n9451), .B(register__n1595), .Y(register__n2794) );
  HB1xp67_ASAP7_75t_R register___U6599 ( .A(register__n8260), .Y(register__n4552) );
  HB1xp67_ASAP7_75t_R register___U6600 ( .A(register__n7928), .Y(register__n5588) );
  INVxp67_ASAP7_75t_R register___U6601 ( .A(register__n1968), .Y(register__n2807) );
  INVxp67_ASAP7_75t_R register___U6602 ( .A(register__n2805), .Y(register__n2817) );
  INVxp33_ASAP7_75t_R register___U6603 ( .A(register__n1957), .Y(register__n2818) );
  INVxp67_ASAP7_75t_R register___U6604 ( .A(register__n2808), .Y(register__n2820) );
  INVxp67_ASAP7_75t_R register___U6605 ( .A(register__n2808), .Y(register__n2821) );
  HB1xp67_ASAP7_75t_R register___U6606 ( .A(register__n2983), .Y(register__n11885) );
  HB1xp67_ASAP7_75t_R register___U6607 ( .A(register__n4587), .Y(register__n2982) );
  HB1xp67_ASAP7_75t_R register___U6608 ( .A(register__n2982), .Y(register__n11884) );
  INVx4_ASAP7_75t_R register___U6609 ( .A(register__n4282), .Y(register__n12263) );
  INVx3_ASAP7_75t_R register___U6610 ( .A(register__net63368), .Y(register__net63324) );
  BUFx3_ASAP7_75t_R register___U6611 ( .A(register__n2831), .Y(register__n2830) );
  BUFx2_ASAP7_75t_R register___U6612 ( .A(register__n10536), .Y(register__n2831) );
  BUFx12f_ASAP7_75t_R register___U6613 ( .A(register__n3248), .Y(register__n11776) );
  BUFx12f_ASAP7_75t_R register___U6614 ( .A(register__n3276), .Y(register__n2840) );
  BUFx3_ASAP7_75t_R register___U6615 ( .A(register__n2842), .Y(register__n2841) );
  BUFx2_ASAP7_75t_R register___U6616 ( .A(register__n11445), .Y(register__n2842) );
  BUFx12f_ASAP7_75t_R register___U6617 ( .A(register__n11781), .Y(register__n2844) );
  BUFx12f_ASAP7_75t_R register___U6618 ( .A(register__n11799), .Y(register__n2846) );
  BUFx3_ASAP7_75t_R register___U6619 ( .A(register__n2848), .Y(register__n2847) );
  BUFx2_ASAP7_75t_R register___U6620 ( .A(register__n11276), .Y(register__n2848) );
  BUFx3_ASAP7_75t_R register___U6621 ( .A(register__n2850), .Y(register__n2849) );
  BUFx2_ASAP7_75t_R register___U6622 ( .A(register__n10939), .Y(register__n2850) );
  BUFx3_ASAP7_75t_R register___U6623 ( .A(register__n2853), .Y(register__n2852) );
  BUFx2_ASAP7_75t_R register___U6624 ( .A(register__n10872), .Y(register__n2853) );
  BUFx12f_ASAP7_75t_R register___U6625 ( .A(register__n11879), .Y(register__n2854) );
  BUFx12f_ASAP7_75t_R register___U6626 ( .A(register__net91920), .Y(register__net64970) );
  INVx6_ASAP7_75t_R register___U6627 ( .A(register__net64870), .Y(register__net64838) );
  BUFx3_ASAP7_75t_R register___U6628 ( .A(register__n2858), .Y(register__n2857) );
  BUFx2_ASAP7_75t_R register___U6629 ( .A(register__n10962), .Y(register__n2858) );
  BUFx3_ASAP7_75t_R register___U6630 ( .A(register__n2861), .Y(register__n2860) );
  BUFx2_ASAP7_75t_R register___U6631 ( .A(register__n10558), .Y(register__n2861) );
  INVx3_ASAP7_75t_R register___U6632 ( .A(register__net64794), .Y(register__net64762) );
  INVx3_ASAP7_75t_R register___U6633 ( .A(register__n12329), .Y(register__n12314) );
  BUFx6f_ASAP7_75t_R register___U6634 ( .A(register__n4639), .Y(register__n12157) );
  INVx6_ASAP7_75t_R register___U6635 ( .A(register__net64452), .Y(register__net64420) );
  INVx6_ASAP7_75t_R register___U6636 ( .A(register__net144463), .Y(register__net64756) );
  INVx6_ASAP7_75t_R register___U6637 ( .A(register__n3259), .Y(register__n11953) );
  INVx6_ASAP7_75t_R register___U6638 ( .A(register__net64036), .Y(register__net64006) );
  INVx6_ASAP7_75t_R register___U6639 ( .A(register__n12300), .Y(register__n12286) );
  BUFx3_ASAP7_75t_R register___U6640 ( .A(register__n2866), .Y(register__n2865) );
  BUFx2_ASAP7_75t_R register___U6641 ( .A(register__n10722), .Y(register__n2866) );
  BUFx3_ASAP7_75t_R register___U6642 ( .A(register__n2868), .Y(register__n2867) );
  BUFx2_ASAP7_75t_R register___U6643 ( .A(register__n11470), .Y(register__n2868) );
  BUFx3_ASAP7_75t_R register___U6644 ( .A(register__n2870), .Y(register__n2869) );
  BUFx2_ASAP7_75t_R register___U6645 ( .A(register__n10768), .Y(register__n2870) );
  INVx6_ASAP7_75t_R register___U6646 ( .A(register__net63220), .Y(register__net63160) );
  INVx3_ASAP7_75t_R register___U6647 ( .A(register__n12215), .Y(register__n12199) );
  INVx3_ASAP7_75t_R register___U6648 ( .A(register__net64764), .Y(register__net147310) );
  BUFx2_ASAP7_75t_R register___U6649 ( .A(register__n2880), .Y(register__n2879) );
  BUFx2_ASAP7_75t_R register___U6650 ( .A(register__n12959), .Y(register__n2880) );
  INVx4_ASAP7_75t_R register___U6651 ( .A(register__n12329), .Y(register__n12317) );
  BUFx12f_ASAP7_75t_R register___U6652 ( .A(register__n2882), .Y(register__n2881) );
  BUFx12f_ASAP7_75t_R register___U6653 ( .A(register__n3277), .Y(register__n2882) );
  INVx3_ASAP7_75t_R register___U6654 ( .A(register__n12408), .Y(register__n12394) );
  BUFx2_ASAP7_75t_R register___U6655 ( .A(register__n10686), .Y(register__n2883) );
  BUFx2_ASAP7_75t_R register___U6656 ( .A(register__n11110), .Y(register__n2887) );
  BUFx2_ASAP7_75t_R register___U6657 ( .A(register__n3409), .Y(register__n2888) );
  BUFx3_ASAP7_75t_R register___U6658 ( .A(register__n2896), .Y(register__n2895) );
  BUFx2_ASAP7_75t_R register___U6659 ( .A(register__n11384), .Y(register__n2896) );
  INVx6_ASAP7_75t_R register___U6660 ( .A(register__net64460), .Y(register__net64416) );
  INVx6_ASAP7_75t_R register___U6661 ( .A(register__net143363), .Y(register__net64836) );
  BUFx2_ASAP7_75t_R register___U6662 ( .A(register__n4038), .Y(register__n2900) );
  INVx6_ASAP7_75t_R register___U6663 ( .A(register__n12268), .Y(register__n12251) );
  BUFx3_ASAP7_75t_R register___U6664 ( .A(register__n2902), .Y(register__n2901) );
  BUFx2_ASAP7_75t_R register___U6665 ( .A(register__n11172), .Y(register__n2902) );
  BUFx2_ASAP7_75t_R register___U6666 ( .A(register__n5538), .Y(register__n2903) );
  BUFx12f_ASAP7_75t_R register___U6667 ( .A(register__net130835), .Y(register__net148409) );
  BUFx3_ASAP7_75t_R register___U6668 ( .A(register__n2905), .Y(register__n2904) );
  BUFx2_ASAP7_75t_R register___U6669 ( .A(register__n11217), .Y(register__n2905) );
  BUFx2_ASAP7_75t_R register___U6670 ( .A(register__n4123), .Y(register__n2906) );
  INVx3_ASAP7_75t_R register___U6671 ( .A(register__n12005), .Y(register__n11989) );
  INVx3_ASAP7_75t_R register___U6672 ( .A(register__n12409), .Y(register__n12399) );
  BUFx3_ASAP7_75t_R register___U6673 ( .A(register__n2910), .Y(register__n2909) );
  BUFx2_ASAP7_75t_R register___U6674 ( .A(register__n11295), .Y(register__n2910) );
  BUFx2_ASAP7_75t_R register___U6675 ( .A(register__n2912), .Y(register__n2911) );
  BUFx2_ASAP7_75t_R register___U6676 ( .A(register__n12898), .Y(register__n2912) );
  BUFx2_ASAP7_75t_R register___U6677 ( .A(register__n2914), .Y(register__n2913) );
  BUFx2_ASAP7_75t_R register___U6678 ( .A(register__n13143), .Y(register__n2914) );
  BUFx2_ASAP7_75t_R register___U6679 ( .A(register__n2916), .Y(register__n2915) );
  BUFx2_ASAP7_75t_R register___U6680 ( .A(register__n12974), .Y(register__n2916) );
  BUFx3_ASAP7_75t_R register___U6681 ( .A(register__n2918), .Y(register__n2917) );
  BUFx2_ASAP7_75t_R register___U6682 ( .A(register__n10983), .Y(register__n2918) );
  BUFx2_ASAP7_75t_R register___U6683 ( .A(register__n2922), .Y(register__n2921) );
  BUFx12f_ASAP7_75t_R register___U6684 ( .A(register__net64052), .Y(register__net64036) );
  BUFx2_ASAP7_75t_R register___U6685 ( .A(register__n2926), .Y(register__n2925) );
  BUFx2_ASAP7_75t_R register___U6686 ( .A(register__n12901), .Y(register__n2926) );
  INVx3_ASAP7_75t_R register___U6687 ( .A(register__n12361), .Y(register__n12349) );
  NOR2x1p5_ASAP7_75t_R register___U6688 ( .A(register__net64430), .B(register__n2813), .Y(register__n8667) );
  BUFx2_ASAP7_75t_R register___U6689 ( .A(register__n2933), .Y(register__n2932) );
  BUFx2_ASAP7_75t_R register___U6690 ( .A(register__n12964), .Y(register__n2933) );
  INVx3_ASAP7_75t_R register___U6691 ( .A(register__net64968), .Y(register__net64934) );
  BUFx2_ASAP7_75t_R register___U6692 ( .A(register__n6263), .Y(register__n2934) );
  BUFx12f_ASAP7_75t_R register___U6693 ( .A(register__n3022), .Y(register__n2935) );
  BUFx2_ASAP7_75t_R register___U6694 ( .A(register__n11067), .Y(register__n2937) );
  BUFx2_ASAP7_75t_R register___U6695 ( .A(register__n3279), .Y(register__n2938) );
  BUFx2_ASAP7_75t_R register___U6696 ( .A(register__n12912), .Y(register__n2940) );
  BUFx2_ASAP7_75t_R register___U6697 ( .A(register__n2942), .Y(register__n2941) );
  BUFx2_ASAP7_75t_R register___U6698 ( .A(register__n2944), .Y(register__n2943) );
  BUFx2_ASAP7_75t_R register___U6699 ( .A(register__n12976), .Y(register__n2944) );
  INVx4_ASAP7_75t_R register___U6700 ( .A(register__n12025), .Y(register__n3501) );
  INVx3_ASAP7_75t_R register___U6701 ( .A(register__n12100), .Y(register__n12087) );
  BUFx2_ASAP7_75t_R register___U6702 ( .A(register__n11023), .Y(register__n2946) );
  BUFx12f_ASAP7_75t_R register___U6703 ( .A(register__n9406), .Y(register__n11970) );
  BUFx2_ASAP7_75t_R register___U6704 ( .A(register__n4472), .Y(register__n2952) );
  INVx6_ASAP7_75t_R register___U6705 ( .A(register__net64384), .Y(register__net64350) );
  INVx3_ASAP7_75t_R register___U6706 ( .A(register__n12103), .Y(register__n12090) );
  BUFx2_ASAP7_75t_R register___U6707 ( .A(register__n11086), .Y(register__n2953) );
  BUFx2_ASAP7_75t_R register___U6708 ( .A(register__n2955), .Y(register__n2954) );
  BUFx2_ASAP7_75t_R register___U6709 ( .A(register__n12918), .Y(register__n2955) );
  INVx3_ASAP7_75t_R register___U6710 ( .A(register__n12157), .Y(register__n12146) );
  INVx3_ASAP7_75t_R register___U6711 ( .A(register__n12360), .Y(register__n12346) );
  INVx3_ASAP7_75t_R register___U6712 ( .A(register__n12382), .Y(register__n12368) );
  INVx6_ASAP7_75t_R register___U6713 ( .A(register__net143690), .Y(register__net64354) );
  BUFx12f_ASAP7_75t_R register___U6714 ( .A(register__n3191), .Y(register__n2967) );
  INVx1_ASAP7_75t_R register___U6715 ( .A(register__n12240), .Y(register__n12228) );
  BUFx2_ASAP7_75t_R register___U6716 ( .A(register__n2974), .Y(register__n2973) );
  BUFx2_ASAP7_75t_R register___U6717 ( .A(register__n12956), .Y(register__n2974) );
  BUFx3_ASAP7_75t_R register___U6718 ( .A(register__n2976), .Y(register__n2975) );
  BUFx2_ASAP7_75t_R register___U6719 ( .A(register__n10538), .Y(register__n2976) );
  BUFx2_ASAP7_75t_R register___U6720 ( .A(register__n7318), .Y(register__n2977) );
  BUFx3_ASAP7_75t_R register___U6721 ( .A(register__n2979), .Y(register__n2978) );
  BUFx2_ASAP7_75t_R register___U6722 ( .A(register__n10537), .Y(register__n2979) );
  BUFx3_ASAP7_75t_R register___U6723 ( .A(register__n2981), .Y(register__n2980) );
  BUFx2_ASAP7_75t_R register___U6724 ( .A(register__n10535), .Y(register__n2981) );
  BUFx2_ASAP7_75t_R register___U6725 ( .A(register__n2990), .Y(register__n2989) );
  BUFx2_ASAP7_75t_R register___U6726 ( .A(register__n13123), .Y(register__n2990) );
  BUFx3_ASAP7_75t_R register___U6727 ( .A(register__n2992), .Y(register__n2991) );
  BUFx2_ASAP7_75t_R register___U6728 ( .A(register__n10829), .Y(register__n2992) );
  BUFx3_ASAP7_75t_R register___U6729 ( .A(register__n2994), .Y(register__n2993) );
  BUFx2_ASAP7_75t_R register___U6730 ( .A(register__n10827), .Y(register__n2994) );
  BUFx3_ASAP7_75t_R register___U6731 ( .A(register__n2996), .Y(register__n2995) );
  BUFx2_ASAP7_75t_R register___U6732 ( .A(register__n10830), .Y(register__n2996) );
  BUFx2_ASAP7_75t_R register___U6733 ( .A(register__n9174), .Y(register__n2997) );
  BUFx3_ASAP7_75t_R register___U6734 ( .A(register__n3001), .Y(register__n3000) );
  BUFx2_ASAP7_75t_R register___U6735 ( .A(register__n11003), .Y(register__n3001) );
  INVx3_ASAP7_75t_R register___U6736 ( .A(register__net63370), .Y(register__net63336) );
  INVx3_ASAP7_75t_R register___U6737 ( .A(register__net63018), .Y(register__net62984) );
  BUFx12f_ASAP7_75t_R register___U6738 ( .A(register__n3542), .Y(register__n3002) );
  BUFx12f_ASAP7_75t_R register___U6739 ( .A(register__n3023), .Y(register__n3003) );
  BUFx12f_ASAP7_75t_R register___U6740 ( .A(register__n3025), .Y(register__n3005) );
  INVx6_ASAP7_75t_R register___U6741 ( .A(register__net63042), .Y(register__net63012) );
  BUFx3_ASAP7_75t_R register___U6742 ( .A(register__n3009), .Y(register__n3008) );
  BUFx2_ASAP7_75t_R register___U6743 ( .A(register__n10724), .Y(register__n3009) );
  BUFx3_ASAP7_75t_R register___U6744 ( .A(register__n3013), .Y(register__n3012) );
  BUFx2_ASAP7_75t_R register___U6745 ( .A(register__n10723), .Y(register__n3013) );
  BUFx3_ASAP7_75t_R register___U6746 ( .A(register__n3015), .Y(register__n3014) );
  BUFx2_ASAP7_75t_R register___U6747 ( .A(register__n10704), .Y(register__n3015) );
  BUFx2_ASAP7_75t_R register___U6748 ( .A(register__n10707), .Y(register__n3016) );
  BUFx2_ASAP7_75t_R register___U6749 ( .A(register__n5377), .Y(register__n3017) );
  BUFx3_ASAP7_75t_R register___U6750 ( .A(register__n3019), .Y(register__n3018) );
  BUFx2_ASAP7_75t_R register___U6751 ( .A(register__n10706), .Y(register__n3019) );
  BUFx6f_ASAP7_75t_R register___U6752 ( .A(register__n3320), .Y(register__n12215) );
  INVx6_ASAP7_75t_R register___U6753 ( .A(register__n3315), .Y(register__n12340) );
  BUFx6f_ASAP7_75t_R register___U6754 ( .A(register__net64798), .Y(register__net64764) );
  BUFx12f_ASAP7_75t_R register___U6755 ( .A(register__n3070), .Y(register__n3023) );
  BUFx12f_ASAP7_75t_R register___U6756 ( .A(register__n3005), .Y(register__n3024) );
  INVx6_ASAP7_75t_R register___U6757 ( .A(register__net63202), .Y(register__net63168) );
  INVx6_ASAP7_75t_R register___U6758 ( .A(register__net145036), .Y(register__net62664) );
  BUFx2_ASAP7_75t_R register___U6759 ( .A(register__n12965), .Y(register__n3029) );
  BUFx3_ASAP7_75t_R register___U6760 ( .A(register__n3031), .Y(register__n3030) );
  BUFx2_ASAP7_75t_R register___U6761 ( .A(register__n7634), .Y(register__n3032) );
  BUFx3_ASAP7_75t_R register___U6762 ( .A(register__n3034), .Y(register__n3033) );
  BUFx2_ASAP7_75t_R register___U6763 ( .A(register__n10920), .Y(register__n3034) );
  BUFx3_ASAP7_75t_R register___U6764 ( .A(register__n3036), .Y(register__n3035) );
  BUFx2_ASAP7_75t_R register___U6765 ( .A(register__n10917), .Y(register__n3036) );
  BUFx3_ASAP7_75t_R register___U6766 ( .A(register__n10769), .Y(register__n3039) );
  BUFx3_ASAP7_75t_R register___U6767 ( .A(register__n3041), .Y(register__n3040) );
  BUFx2_ASAP7_75t_R register___U6768 ( .A(register__n10770), .Y(register__n3041) );
  BUFx2_ASAP7_75t_R register___U6769 ( .A(register__n3643), .Y(register__n3042) );
  INVx3_ASAP7_75t_R register___U6770 ( .A(register__n12363), .Y(register__n12348) );
  INVx3_ASAP7_75t_R register___U6771 ( .A(register__n12411), .Y(register__n12400) );
  BUFx12f_ASAP7_75t_R register___U6772 ( .A(register__n3218), .Y(register__n3044) );
  INVx6_ASAP7_75t_R register___U6773 ( .A(register__net146116), .Y(register__net64328) );
  BUFx2_ASAP7_75t_R register___U6774 ( .A(register__n12954), .Y(register__n3045) );
  BUFx2_ASAP7_75t_R register___U6775 ( .A(register__n3563), .Y(register__n3050) );
  BUFx2_ASAP7_75t_R register___U6776 ( .A(register__n12978), .Y(register__n3051) );
  BUFx3_ASAP7_75t_R register___U6777 ( .A(register__n3057), .Y(register__n3056) );
  BUFx2_ASAP7_75t_R register___U6778 ( .A(register__n11537), .Y(register__n3057) );
  BUFx3_ASAP7_75t_R register___U6779 ( .A(register__n3059), .Y(register__n3058) );
  BUFx2_ASAP7_75t_R register___U6780 ( .A(register__n10848), .Y(register__n3059) );
  BUFx3_ASAP7_75t_R register___U6781 ( .A(register__n3062), .Y(register__n3061) );
  BUFx2_ASAP7_75t_R register___U6782 ( .A(register__n10850), .Y(register__n3062) );
  BUFx3_ASAP7_75t_R register___U6783 ( .A(register__n3065), .Y(register__n3064) );
  BUFx2_ASAP7_75t_R register___U6784 ( .A(register__n10984), .Y(register__n3065) );
  BUFx3_ASAP7_75t_R register___U6785 ( .A(register__n3067), .Y(register__n3066) );
  BUFx2_ASAP7_75t_R register___U6786 ( .A(register__n10982), .Y(register__n3067) );
  BUFx12f_ASAP7_75t_R register___U6787 ( .A(register__n3003), .Y(register__n3068) );
  INVx6_ASAP7_75t_R register___U6788 ( .A(register__net64368), .Y(register__net64336) );
  BUFx12f_ASAP7_75t_R register___U6789 ( .A(register__net117320), .Y(register__net64368) );
  INVx3_ASAP7_75t_R register___U6790 ( .A(register__n11977), .Y(register__n11963) );
  INVx6_ASAP7_75t_R register___U6791 ( .A(register__n3314), .Y(register__n12342) );
  INVx5_ASAP7_75t_R register___U6792 ( .A(register__n11970), .Y(register__n11955) );
  INVx6_ASAP7_75t_R register___U6793 ( .A(register__net64030), .Y(register__net64004) );
  BUFx2_ASAP7_75t_R register___U6794 ( .A(register__n4484), .Y(register__n3079) );
  BUFx2_ASAP7_75t_R register___U6795 ( .A(register__n12953), .Y(register__n3080) );
  BUFx2_ASAP7_75t_R register___U6796 ( .A(register__n3751), .Y(register__n3081) );
  BUFx2_ASAP7_75t_R register___U6797 ( .A(register__n5238), .Y(register__n3082) );
  BUFx2_ASAP7_75t_R register___U6798 ( .A(register__n12975), .Y(register__n3083) );
  BUFx3_ASAP7_75t_R register___U6799 ( .A(register__n3085), .Y(register__n3084) );
  BUFx2_ASAP7_75t_R register___U6800 ( .A(register__n11491), .Y(register__n3085) );
  BUFx3_ASAP7_75t_R register___U6801 ( .A(register__n3087), .Y(register__n3086) );
  BUFx2_ASAP7_75t_R register___U6802 ( .A(register__n11493), .Y(register__n3087) );
  BUFx2_ASAP7_75t_R register___U6803 ( .A(register__n7636), .Y(register__n3088) );
  BUFx3_ASAP7_75t_R register___U6804 ( .A(register__n3090), .Y(register__n3089) );
  BUFx2_ASAP7_75t_R register___U6805 ( .A(register__n11490), .Y(register__n3090) );
  BUFx3_ASAP7_75t_R register___U6806 ( .A(register__n3092), .Y(register__n3091) );
  BUFx2_ASAP7_75t_R register___U6807 ( .A(register__n10873), .Y(register__n3092) );
  BUFx3_ASAP7_75t_R register___U6808 ( .A(register__n3096), .Y(register__n3095) );
  BUFx2_ASAP7_75t_R register___U6809 ( .A(register__n10871), .Y(register__n3096) );
  BUFx3_ASAP7_75t_R register___U6810 ( .A(register__n3098), .Y(register__n3097) );
  BUFx2_ASAP7_75t_R register___U6811 ( .A(register__n10964), .Y(register__n3098) );
  BUFx3_ASAP7_75t_R register___U6812 ( .A(register__n3100), .Y(register__n3099) );
  BUFx2_ASAP7_75t_R register___U6813 ( .A(register__n10963), .Y(register__n3100) );
  BUFx3_ASAP7_75t_R register___U6814 ( .A(register__n3102), .Y(register__n3101) );
  BUFx2_ASAP7_75t_R register___U6815 ( .A(register__n10961), .Y(register__n3102) );
  BUFx2_ASAP7_75t_R register___U6816 ( .A(register__n10688), .Y(register__n3103) );
  BUFx3_ASAP7_75t_R register___U6817 ( .A(register__n3105), .Y(register__n3104) );
  BUFx2_ASAP7_75t_R register___U6818 ( .A(register__n10687), .Y(register__n3105) );
  BUFx2_ASAP7_75t_R register___U6819 ( .A(register__n11024), .Y(register__n3108) );
  BUFx3_ASAP7_75t_R register___U6820 ( .A(register__n3113), .Y(register__n3112) );
  BUFx2_ASAP7_75t_R register___U6821 ( .A(register__n11654), .Y(register__n3113) );
  BUFx3_ASAP7_75t_R register___U6822 ( .A(register__n3115), .Y(register__n3114) );
  BUFx2_ASAP7_75t_R register___U6823 ( .A(register__n11696), .Y(register__n3115) );
  INVx3_ASAP7_75t_R register___U6824 ( .A(register__n11976), .Y(register__n11960) );
  BUFx12f_ASAP7_75t_R register___U6825 ( .A(register__net145767), .Y(register__net146677) );
  BUFx3_ASAP7_75t_R register___U6826 ( .A(register__n3122), .Y(register__n3121) );
  BUFx2_ASAP7_75t_R register___U6827 ( .A(register__n10577), .Y(register__n3122) );
  BUFx2_ASAP7_75t_R register___U6828 ( .A(register__n3124), .Y(register__n3123) );
  BUFx2_ASAP7_75t_R register___U6829 ( .A(register__n13132), .Y(register__n3124) );
  BUFx2_ASAP7_75t_R register___U6830 ( .A(register__n10603), .Y(register__n3131) );
  BUFx3_ASAP7_75t_R register___U6831 ( .A(register__n10940), .Y(register__n3132) );
  BUFx3_ASAP7_75t_R register___U6832 ( .A(register__n3134), .Y(register__n3133) );
  BUFx2_ASAP7_75t_R register___U6833 ( .A(register__n10941), .Y(register__n3134) );
  BUFx3_ASAP7_75t_R register___U6834 ( .A(register__n3136), .Y(register__n3135) );
  BUFx2_ASAP7_75t_R register___U6835 ( .A(register__n10938), .Y(register__n3136) );
  BUFx3_ASAP7_75t_R register___U6836 ( .A(register__n3138), .Y(register__n3137) );
  BUFx2_ASAP7_75t_R register___U6837 ( .A(register__n10896), .Y(register__n3138) );
  BUFx3_ASAP7_75t_R register___U6838 ( .A(register__n3140), .Y(register__n3139) );
  BUFx2_ASAP7_75t_R register___U6839 ( .A(register__n10894), .Y(register__n3140) );
  BUFx2_ASAP7_75t_R register___U6840 ( .A(register__n11427), .Y(register__n3143) );
  BUFx3_ASAP7_75t_R register___U6841 ( .A(register__n3145), .Y(register__n3144) );
  BUFx2_ASAP7_75t_R register___U6842 ( .A(register__n11085), .Y(register__n3145) );
  BUFx2_ASAP7_75t_R register___U6843 ( .A(register__n11087), .Y(register__n3146) );
  BUFx12f_ASAP7_75t_R register___U6844 ( .A(register__n2985), .Y(register__n3148) );
  BUFx12f_ASAP7_75t_R register___U6845 ( .A(register__n3150), .Y(register__n3149) );
  BUFx12f_ASAP7_75t_R register___U6846 ( .A(register__n4031), .Y(register__n3150) );
  BUFx12f_ASAP7_75t_R register___U6847 ( .A(register__n3219), .Y(register__n4031) );
  INVx3_ASAP7_75t_R register___U6848 ( .A(register__net64386), .Y(register__net64356) );
  BUFx12f_ASAP7_75t_R register___U6849 ( .A(register__n3155), .Y(register__n3154) );
  BUFx12f_ASAP7_75t_R register___U6850 ( .A(register__n3192), .Y(register__n3155) );
  BUFx2_ASAP7_75t_R register___U6851 ( .A(register__n3161), .Y(register__n3160) );
  BUFx2_ASAP7_75t_R register___U6852 ( .A(register__n13364), .Y(register__n3161) );
  CKINVDCx10_ASAP7_75t_R register___U6853 ( .A(register__net63214), .Y(register__net63178) );
  BUFx2_ASAP7_75t_R register___U6854 ( .A(register__n10918), .Y(register__n3166) );
  BUFx2_ASAP7_75t_R register___U6855 ( .A(register__n8275), .Y(register__n3167) );
  BUFx4f_ASAP7_75t_R register___U6856 ( .A(register__net63330), .Y(register__net146308) );
  BUFx12f_ASAP7_75t_R register___U6857 ( .A(register__net146408), .Y(register__net146266) );
  BUFx12f_ASAP7_75t_R register___U6858 ( .A(register__net146266), .Y(register__net64460) );
  BUFx2_ASAP7_75t_R register___U6859 ( .A(register__n3173), .Y(register__n3172) );
  BUFx2_ASAP7_75t_R register___U6860 ( .A(register__n13367), .Y(register__n3173) );
  BUFx2_ASAP7_75t_R register___U6861 ( .A(register__n3176), .Y(register__n3175) );
  BUFx2_ASAP7_75t_R register___U6862 ( .A(register__n13128), .Y(register__n3176) );
  BUFx2_ASAP7_75t_R register___U6863 ( .A(register__n11723), .Y(register__n3179) );
  BUFx2_ASAP7_75t_R register___U6864 ( .A(register__n11722), .Y(register__n3181) );
  INVx2_ASAP7_75t_R register___U6865 ( .A(register__n3475), .Y(register__n3186) );
  INVx6_ASAP7_75t_R register___U6866 ( .A(register__net64876), .Y(register__net64844) );
  BUFx12f_ASAP7_75t_R register___U6867 ( .A(register__net64378), .Y(register__net146116) );
  BUFx12f_ASAP7_75t_R register___U6868 ( .A(register__n2962), .Y(register__n3188) );
  BUFx12f_ASAP7_75t_R register___U6869 ( .A(register__n3157), .Y(register__n11968) );
  BUFx12f_ASAP7_75t_R register___U6870 ( .A(register__n11850), .Y(register__n3191) );
  BUFx12f_ASAP7_75t_R register___U6871 ( .A(register__n3316), .Y(register__n3192) );
  BUFx2_ASAP7_75t_R register___U6872 ( .A(register__n3194), .Y(register__n3193) );
  BUFx2_ASAP7_75t_R register___U6873 ( .A(register__n12810), .Y(register__n3194) );
  BUFx2_ASAP7_75t_R register___U6874 ( .A(register__n3198), .Y(register__n3197) );
  BUFx2_ASAP7_75t_R register___U6875 ( .A(register__n13137), .Y(register__n3198) );
  BUFx3_ASAP7_75t_R register___U6876 ( .A(register__n3201), .Y(register__n3200) );
  BUFx2_ASAP7_75t_R register___U6877 ( .A(register__n11579), .Y(register__n3201) );
  BUFx2_ASAP7_75t_R register___U6878 ( .A(register__n5695), .Y(register__n3202) );
  BUFx3_ASAP7_75t_R register___U6879 ( .A(register__n3204), .Y(register__n3203) );
  BUFx2_ASAP7_75t_R register___U6880 ( .A(register__n11577), .Y(register__n3204) );
  BUFx3_ASAP7_75t_R register___U6881 ( .A(register__n3206), .Y(register__n3205) );
  BUFx2_ASAP7_75t_R register___U6882 ( .A(register__n11446), .Y(register__n3206) );
  BUFx3_ASAP7_75t_R register___U6883 ( .A(register__n3208), .Y(register__n3207) );
  BUFx3_ASAP7_75t_R register___U6884 ( .A(register__n8166), .Y(register__n3213) );
  BUFx6f_ASAP7_75t_R register___U6885 ( .A(register__n8165), .Y(register__n9842) );
  BUFx4f_ASAP7_75t_R register___U6886 ( .A(register__n3213), .Y(register__n8165) );
  BUFx6f_ASAP7_75t_R register___U6887 ( .A(register__net64804), .Y(register__net127692) );
  BUFx3_ASAP7_75t_R register___U6888 ( .A(register__n3841), .Y(register__n3214) );
  BUFx3_ASAP7_75t_R register___U6889 ( .A(register__n3841), .Y(register__n3215) );
  INVx3_ASAP7_75t_R register___U6890 ( .A(register__n12358), .Y(register__n12345) );
  BUFx12f_ASAP7_75t_R register___U6891 ( .A(register__n3189), .Y(register__n3218) );
  BUFx12f_ASAP7_75t_R register___U6892 ( .A(register__net100540), .Y(register__net145767) );
  BUFx2_ASAP7_75t_R register___U6893 ( .A(register__n3223), .Y(register__n3222) );
  BUFx2_ASAP7_75t_R register___U6894 ( .A(register__n13371), .Y(register__n3223) );
  BUFx2_ASAP7_75t_R register___U6895 ( .A(register__n3225), .Y(register__n3224) );
  BUFx2_ASAP7_75t_R register___U6896 ( .A(register__n12900), .Y(register__n3225) );
  BUFx2_ASAP7_75t_R register___U6897 ( .A(register__n3227), .Y(register__n3226) );
  BUFx2_ASAP7_75t_R register___U6898 ( .A(register__n13124), .Y(register__n3227) );
  BUFx3_ASAP7_75t_R register___U6899 ( .A(register__n3231), .Y(register__n3230) );
  BUFx2_ASAP7_75t_R register___U6900 ( .A(register__n11194), .Y(register__n3231) );
  BUFx3_ASAP7_75t_R register___U6901 ( .A(register__n3233), .Y(register__n3232) );
  BUFx2_ASAP7_75t_R register___U6902 ( .A(register__n11192), .Y(register__n3233) );
  BUFx2_ASAP7_75t_R register___U6903 ( .A(register__n11382), .Y(register__n3244) );
  BUFx2_ASAP7_75t_R register___U6904 ( .A(register__n8227), .Y(register__n3247) );
  BUFx12f_ASAP7_75t_R register___U6905 ( .A(register__n11878), .Y(register__n3248) );
  BUFx12f_ASAP7_75t_R register___U6906 ( .A(register__n11880), .Y(register__n11878) );
  BUFx3_ASAP7_75t_R register___U6907 ( .A(register__n7764), .Y(register__n3249) );
  BUFx6f_ASAP7_75t_R register___U6908 ( .A(register__n7763), .Y(register__n10003) );
  BUFx4f_ASAP7_75t_R register___U6909 ( .A(register__n3249), .Y(register__n7763) );
  BUFx3_ASAP7_75t_R register___U6910 ( .A(register__n7812), .Y(register__n3250) );
  BUFx4f_ASAP7_75t_R register___U6911 ( .A(register__n3250), .Y(register__n7811) );
  BUFx3_ASAP7_75t_R register___U6912 ( .A(register__n5215), .Y(register__n3251) );
  BUFx3_ASAP7_75t_R register___U6913 ( .A(register__n8545), .Y(register__n3252) );
  BUFx6f_ASAP7_75t_R register___U6914 ( .A(register__n9902), .Y(register__n9901) );
  BUFx4f_ASAP7_75t_R register___U6915 ( .A(register__n12123), .Y(register__n3253) );
  BUFx12f_ASAP7_75t_R register___U6916 ( .A(register__n12154), .Y(register__n3255) );
  BUFx12f_ASAP7_75t_R register___U6917 ( .A(register__net145772), .Y(register__net145521) );
  BUFx12f_ASAP7_75t_R register___U6918 ( .A(register__net145773), .Y(register__net145522) );
  BUFx12f_ASAP7_75t_R register___U6919 ( .A(register__net64884), .Y(register__net145523) );
  BUFx12f_ASAP7_75t_R register___U6920 ( .A(register__net145521), .Y(register__net64876) );
  INVx3_ASAP7_75t_R register___U6921 ( .A(register__n12479), .Y(register__n12463) );
  BUFx12f_ASAP7_75t_R register___U6922 ( .A(register__n11969), .Y(register__n3260) );
  BUFx12f_ASAP7_75t_R register___U6923 ( .A(register__n3282), .Y(register__n3262) );
  BUFx12f_ASAP7_75t_R register___U6924 ( .A(register__n8334), .Y(register__n3879) );
  BUFx12f_ASAP7_75t_R register___U6925 ( .A(register__n11814), .Y(register__n3268) );
  BUFx2_ASAP7_75t_R register___U6926 ( .A(register__n3270), .Y(register__n3269) );
  BUFx2_ASAP7_75t_R register___U6927 ( .A(register__n13381), .Y(register__n3270) );
  BUFx12f_ASAP7_75t_R register___U6928 ( .A(register__n12391), .Y(register__n3273) );
  BUFx12f_ASAP7_75t_R register___U6929 ( .A(register__n3273), .Y(register__n12384) );
  BUFx12f_ASAP7_75t_R register___U6930 ( .A(register__n2840), .Y(register__n3274) );
  BUFx12f_ASAP7_75t_R register___U6931 ( .A(register__n11779), .Y(register__n11778) );
  BUFx12f_ASAP7_75t_R register___U6932 ( .A(register__n11778), .Y(register__n11879) );
  INVx1_ASAP7_75t_R register___U6933 ( .A(register__n2937), .Y(register__n3279) );
  INVx3_ASAP7_75t_R register___U6934 ( .A(register__n12129), .Y(register__n12113) );
  BUFx12f_ASAP7_75t_R register___U6935 ( .A(register__net129615), .Y(register__net62682) );
  INVx3_ASAP7_75t_R register___U6936 ( .A(register__net63380), .Y(register__net63344) );
  INVx6_ASAP7_75t_R register___U6937 ( .A(register__n12159), .Y(register__n12148) );
  BUFx12f_ASAP7_75t_R register___U6938 ( .A(register__n3148), .Y(register__n12159) );
  BUFx12f_ASAP7_75t_R register___U6939 ( .A(register__net145247), .Y(register__net145245) );
  BUFx12f_ASAP7_75t_R register___U6940 ( .A(register__net64896), .Y(register__net145247) );
  BUFx12f_ASAP7_75t_R register___U6941 ( .A(register__n12476), .Y(register__n3281) );
  BUFx12f_ASAP7_75t_R register___U6942 ( .A(register__n3708), .Y(register__n3282) );
  BUFx12f_ASAP7_75t_R register___U6943 ( .A(register__n3545), .Y(register__n3284) );
  BUFx12f_ASAP7_75t_R register___U6944 ( .A(register__net145449), .Y(register__net145201) );
  BUFx12f_ASAP7_75t_R register___U6945 ( .A(register__net144689), .Y(register__net145202) );
  BUFx2_ASAP7_75t_R register___U6946 ( .A(register__n3288), .Y(register__n3287) );
  BUFx2_ASAP7_75t_R register___U6947 ( .A(register__n12823), .Y(register__n3288) );
  BUFx2_ASAP7_75t_R register___U6948 ( .A(register__n3290), .Y(register__n3289) );
  BUFx2_ASAP7_75t_R register___U6949 ( .A(register__n13001), .Y(register__n3290) );
  BUFx2_ASAP7_75t_R register___U6950 ( .A(register__n3292), .Y(register__n3291) );
  BUFx2_ASAP7_75t_R register___U6951 ( .A(register__n13383), .Y(register__n3292) );
  INVx1_ASAP7_75t_R register___U6952 ( .A(register__n2852), .Y(register__n3303) );
  BUFx6f_ASAP7_75t_R register___U6953 ( .A(register__n4650), .Y(register__n12209) );
  INVx3_ASAP7_75t_R register___U6954 ( .A(register__net64054), .Y(register__net64018) );
  BUFx6f_ASAP7_75t_R register___U6955 ( .A(register__net64038), .Y(register__net64054) );
  INVx2_ASAP7_75t_R register___U6956 ( .A(register__n3838), .Y(register__n3305) );
  INVx6_ASAP7_75t_R register___U6957 ( .A(register__n3629), .Y(register__n12110) );
  BUFx12f_ASAP7_75t_R register___U6958 ( .A(register__net145038), .Y(register__net145036) );
  BUFx12f_ASAP7_75t_R register___U6959 ( .A(register__net145038), .Y(register__net145037) );
  BUFx12f_ASAP7_75t_R register___U6960 ( .A(register__net62698), .Y(register__net145038) );
  INVx3_ASAP7_75t_R register___U6961 ( .A(register__net63270), .Y(register__net63236) );
  INVx3_ASAP7_75t_R register___U6962 ( .A(register__n12296), .Y(register__n12282) );
  BUFx12f_ASAP7_75t_R register___U6963 ( .A(register__n3281), .Y(register__n4000) );
  INVx6_ASAP7_75t_R register___U6964 ( .A(register__net64954), .Y(register__net64922) );
  BUFx12f_ASAP7_75t_R register___U6965 ( .A(register__net91923), .Y(register__net64954) );
  BUFx12f_ASAP7_75t_R register___U6966 ( .A(register__net144717), .Y(register__net144981) );
  INVx6_ASAP7_75t_R register___U6967 ( .A(register__n3356), .Y(register__n12281) );
  BUFx12f_ASAP7_75t_R register___U6968 ( .A(register__net142573), .Y(register__net142960) );
  BUFx2_ASAP7_75t_R register___U6969 ( .A(register__n3311), .Y(register__n3310) );
  BUFx2_ASAP7_75t_R register___U6970 ( .A(register__n12731), .Y(register__n3311) );
  BUFx2_ASAP7_75t_R register___U6971 ( .A(register__n3313), .Y(register__n3312) );
  BUFx2_ASAP7_75t_R register___U6972 ( .A(register__n12825), .Y(register__n3313) );
  BUFx12f_ASAP7_75t_R register___U6973 ( .A(register__n3266), .Y(register__n3314) );
  BUFx12f_ASAP7_75t_R register___U6974 ( .A(register__n12354), .Y(register__n3315) );
  BUFx12f_ASAP7_75t_R register___U6975 ( .A(register__n3317), .Y(register__n11880) );
  INVx1_ASAP7_75t_R register___U6976 ( .A(register__n2857), .Y(register__n3318) );
  BUFx4f_ASAP7_75t_R register___U6977 ( .A(register__n12423), .Y(register__n3319) );
  BUFx12f_ASAP7_75t_R register___U6978 ( .A(register__n12305), .Y(register__n3321) );
  BUFx12f_ASAP7_75t_R register___U6979 ( .A(register__n12305), .Y(register__n3322) );
  INVx4_ASAP7_75t_R register___U6980 ( .A(register__n3321), .Y(register__n12279) );
  INVx3_ASAP7_75t_R register___U6981 ( .A(register__n12270), .Y(register__n12257) );
  INVx3_ASAP7_75t_R register___U6982 ( .A(register__n12186), .Y(register__n12174) );
  BUFx12f_ASAP7_75t_R register___U6983 ( .A(register__n12481), .Y(register__n3323) );
  INVx2_ASAP7_75t_R register___U6984 ( .A(register__n3323), .Y(register__n12465) );
  BUFx4f_ASAP7_75t_R register___U6985 ( .A(register__n12481), .Y(register__n12466) );
  BUFx12f_ASAP7_75t_R register___U6986 ( .A(register__n11763), .Y(register__n3324) );
  BUFx12f_ASAP7_75t_R register___U6987 ( .A(register__n5342), .Y(register__n3325) );
  BUFx12f_ASAP7_75t_R register___U6988 ( .A(register__net141026), .Y(register__net144717) );
  BUFx12f_ASAP7_75t_R register___U6989 ( .A(register__net145246), .Y(register__net102923) );
  BUFx2_ASAP7_75t_R register___U6990 ( .A(register__n3331), .Y(register__n3330) );
  INVx6_ASAP7_75t_R register___U6991 ( .A(register__net64882), .Y(register__net64848) );
  BUFx12f_ASAP7_75t_R register___U6992 ( .A(register__net136187), .Y(register__net144561) );
  BUFx12f_ASAP7_75t_R register___U6993 ( .A(register__net136187), .Y(register__net144562) );
  BUFx12f_ASAP7_75t_R register___U6994 ( .A(register__net144562), .Y(register__net63024) );
  BUFx12f_ASAP7_75t_R register___U6995 ( .A(register__n3154), .Y(register__n3341) );
  INVx1_ASAP7_75t_R register___U6996 ( .A(register__n2893), .Y(register__n3345) );
  INVx6_ASAP7_75t_R register___U6997 ( .A(register__net143695), .Y(register__net63996) );
  INVx4_ASAP7_75t_R register___U6998 ( .A(register__net141387), .Y(register__net63014) );
  INVx3_ASAP7_75t_R register___U6999 ( .A(register__n12328), .Y(register__n12316) );
  INVx3_ASAP7_75t_R register___U7000 ( .A(register__n12007), .Y(register__n11985) );
  INVx3_ASAP7_75t_R register___U7001 ( .A(register__n12442), .Y(register__n12426) );
  BUFx12f_ASAP7_75t_R register___U7002 ( .A(register__n12355), .Y(register__n3347) );
  INVx2_ASAP7_75t_R register___U7003 ( .A(register__n3346), .Y(register__n4999) );
  BUFx12f_ASAP7_75t_R register___U7004 ( .A(register__n6430), .Y(register__n3351) );
  BUFx12f_ASAP7_75t_R register___U7005 ( .A(register__n3357), .Y(register__n3355) );
  BUFx12f_ASAP7_75t_R register___U7006 ( .A(register__n3358), .Y(register__n3356) );
  BUFx12f_ASAP7_75t_R register___U7007 ( .A(register__n3361), .Y(register__n3360) );
  BUFx12f_ASAP7_75t_R register___U7008 ( .A(register__n11843), .Y(register__n3361) );
  BUFx12f_ASAP7_75t_R register___U7009 ( .A(register__n3427), .Y(register__n3362) );
  BUFx12f_ASAP7_75t_R register___U7010 ( .A(register__n3379), .Y(register__n3366) );
  INVx6_ASAP7_75t_R register___U7011 ( .A(register__n12067), .Y(register__n12053) );
  INVx5_ASAP7_75t_R register___U7012 ( .A(register__net64372), .Y(register__net64340) );
  BUFx2_ASAP7_75t_R register___U7013 ( .A(register__n3370), .Y(register__n3369) );
  BUFx2_ASAP7_75t_R register___U7014 ( .A(register__n13365), .Y(register__n3370) );
  INVx1_ASAP7_75t_R register___U7015 ( .A(register__n3121), .Y(register__n3372) );
  BUFx12f_ASAP7_75t_R register___U7016 ( .A(register__n708), .Y(register__n11779) );
  INVx4_ASAP7_75t_R register___U7017 ( .A(register__n108), .Y(register__n12176) );
  BUFx12f_ASAP7_75t_R register___U7018 ( .A(register__n3365), .Y(register__n3377) );
  INVx4_ASAP7_75t_R register___U7019 ( .A(register__n12302), .Y(register__n12287) );
  INVx3_ASAP7_75t_R register___U7020 ( .A(register__n12443), .Y(register__n12427) );
  INVx3_ASAP7_75t_R register___U7021 ( .A(register__net63374), .Y(register__net63340) );
  INVx2_ASAP7_75t_R register___U7022 ( .A(register__n12467), .Y(register__n12451) );
  BUFx12f_ASAP7_75t_R register___U7023 ( .A(register__net144158), .Y(register__net144157) );
  BUFx12f_ASAP7_75t_R register___U7024 ( .A(register__net136275), .Y(register__net144158) );
  BUFx12f_ASAP7_75t_R register___U7025 ( .A(register__n3680), .Y(register__n3382) );
  BUFx12f_ASAP7_75t_R register___U7026 ( .A(register__n3421), .Y(register__n3386) );
  BUFx12f_ASAP7_75t_R register___U7027 ( .A(register__n12095), .Y(register__n3387) );
  BUFx6f_ASAP7_75t_R register___U7028 ( .A(register__n12095), .Y(register__n3388) );
  INVx2_ASAP7_75t_R register___U7029 ( .A(register__n3388), .Y(register__n12085) );
  BUFx12f_ASAP7_75t_R register___U7030 ( .A(register__n3254), .Y(register__n4848) );
  BUFx2_ASAP7_75t_R register___U7031 ( .A(register__n3397), .Y(register__n3396) );
  INVx6_ASAP7_75t_R register___U7032 ( .A(register__net63194), .Y(register__net63162) );
  BUFx2_ASAP7_75t_R register___U7033 ( .A(register__n3399), .Y(register__n3398) );
  BUFx2_ASAP7_75t_R register___U7034 ( .A(register__n13005), .Y(register__n3399) );
  INVx4_ASAP7_75t_R register___U7035 ( .A(register__n3323), .Y(register__n12453) );
  BUFx2_ASAP7_75t_R register___U7036 ( .A(register__n3403), .Y(register__n3402) );
  BUFx2_ASAP7_75t_R register___U7037 ( .A(register__n13379), .Y(register__n3403) );
  BUFx2_ASAP7_75t_R register___U7038 ( .A(register__n4980), .Y(register__n3406) );
  INVx6_ASAP7_75t_R register___U7039 ( .A(register__net63200), .Y(register__net63156) );
  BUFx12f_ASAP7_75t_R register___U7040 ( .A(register__n11797), .Y(register__n11883) );
  INVx1_ASAP7_75t_R register___U7041 ( .A(register__n2887), .Y(register__n3409) );
  INVx6_ASAP7_75t_R register___U7042 ( .A(register__n11940), .Y(register__n11923) );
  BUFx12f_ASAP7_75t_R register___U7043 ( .A(register__n11937), .Y(register__n11940) );
  BUFx2_ASAP7_75t_R register___U7044 ( .A(register__n12255), .Y(register__n3411) );
  INVx6_ASAP7_75t_R register___U7045 ( .A(register__n3531), .Y(register__n12406) );
  BUFx12f_ASAP7_75t_R register___U7046 ( .A(register__n7609), .Y(register__n3412) );
  BUFx12f_ASAP7_75t_R register___U7047 ( .A(register__n3412), .Y(register__n11975) );
  BUFx12f_ASAP7_75t_R register___U7048 ( .A(register__net97625), .Y(register__net129770) );
  BUFx12f_ASAP7_75t_R register___U7049 ( .A(register__n5342), .Y(register__n3415) );
  BUFx12f_ASAP7_75t_R register___U7050 ( .A(register__n3417), .Y(register__n3416) );
  BUFx12f_ASAP7_75t_R register___U7051 ( .A(register__n3349), .Y(register__n3417) );
  BUFx12f_ASAP7_75t_R register___U7052 ( .A(register__n3386), .Y(register__n3420) );
  BUFx12f_ASAP7_75t_R register___U7053 ( .A(register__n3517), .Y(register__n3421) );
  BUFx12f_ASAP7_75t_R register___U7054 ( .A(register__net129691), .Y(register__net143813) );
  BUFx12f_ASAP7_75t_R register___U7055 ( .A(register__net143517), .Y(register__net143789) );
  BUFx12f_ASAP7_75t_R register___U7056 ( .A(register__n3450), .Y(register__n3424) );
  BUFx12f_ASAP7_75t_R register___U7057 ( .A(register__n12096), .Y(register__n3427) );
  BUFx12f_ASAP7_75t_R register___U7058 ( .A(register__net74027), .Y(register__net143769) );
  INVx6_ASAP7_75t_R register___U7059 ( .A(register__net62686), .Y(register__net62654) );
  BUFx2_ASAP7_75t_R register___U7060 ( .A(register__n3429), .Y(register__n3428) );
  INVx6_ASAP7_75t_R register___U7061 ( .A(register__net64888), .Y(register__net64854) );
  BUFx2_ASAP7_75t_R register___U7062 ( .A(register__n3435), .Y(register__n3434) );
  BUFx2_ASAP7_75t_R register___U7063 ( .A(register__n13366), .Y(register__n3435) );
  BUFx12f_ASAP7_75t_R register___U7064 ( .A(register__net130835), .Y(register__net143694) );
  BUFx12f_ASAP7_75t_R register___U7065 ( .A(register__net64040), .Y(register__net143695) );
  BUFx12f_ASAP7_75t_R register___U7066 ( .A(register__net64390), .Y(register__net143690) );
  BUFx12f_ASAP7_75t_R register___U7067 ( .A(register__n3274), .Y(register__n11869) );
  BUFx4f_ASAP7_75t_R register___U7068 ( .A(register__n12024), .Y(register__n3441) );
  INVx2_ASAP7_75t_R register___U7069 ( .A(register__n3594), .Y(register__n3442) );
  BUFx12f_ASAP7_75t_R register___U7070 ( .A(register__net144161), .Y(register__net63220) );
  INVx3_ASAP7_75t_R register___U7071 ( .A(register__net64806), .Y(register__net64776) );
  BUFx6f_ASAP7_75t_R register___U7072 ( .A(register__n12179), .Y(register__n12166) );
  INVx3_ASAP7_75t_R register___U7073 ( .A(register__n12166), .Y(register__n3445) );
  INVx3_ASAP7_75t_R register___U7074 ( .A(register__net62872), .Y(register__net62838) );
  BUFx12f_ASAP7_75t_R register___U7075 ( .A(register__n7296), .Y(register__n3447) );
  BUFx12f_ASAP7_75t_R register___U7076 ( .A(register__net143789), .Y(register__net143516) );
  BUFx12f_ASAP7_75t_R register___U7077 ( .A(register__net140597), .Y(register__net143517) );
  BUFx12f_ASAP7_75t_R register___U7078 ( .A(register__n3424), .Y(register__n3448) );
  BUFx12f_ASAP7_75t_R register___U7079 ( .A(register__n12472), .Y(register__n3450) );
  BUFx12f_ASAP7_75t_R register___U7080 ( .A(register__n3473), .Y(register__n3452) );
  BUFx12f_ASAP7_75t_R register___U7081 ( .A(register__net143492), .Y(register__net143491) );
  BUFx12f_ASAP7_75t_R register___U7082 ( .A(register__net139025), .Y(register__net143492) );
  BUFx12f_ASAP7_75t_R register___U7083 ( .A(register__n3483), .Y(register__n3455) );
  BUFx12f_ASAP7_75t_R register___U7084 ( .A(register__n3156), .Y(register__n11971) );
  BUFx2_ASAP7_75t_R register___U7085 ( .A(register__n3459), .Y(register__n3458) );
  BUFx2_ASAP7_75t_R register___U7086 ( .A(register__n3463), .Y(register__n3462) );
  BUFx2_ASAP7_75t_R register___U7087 ( .A(register__n12818), .Y(register__n3463) );
  BUFx2_ASAP7_75t_R register___U7088 ( .A(register__n3465), .Y(register__n3464) );
  BUFx2_ASAP7_75t_R register___U7089 ( .A(register__n13380), .Y(register__n3465) );
  BUFx2_ASAP7_75t_R register___U7090 ( .A(register__n5494), .Y(register__n3468) );
  INVx3_ASAP7_75t_R register___U7091 ( .A(register__net64808), .Y(register__net64772) );
  INVx3_ASAP7_75t_R register___U7092 ( .A(register__net64050), .Y(register__net64020) );
  INVx3_ASAP7_75t_R register___U7093 ( .A(register__n12187), .Y(register__n12177) );
  INVx3_ASAP7_75t_R register___U7094 ( .A(register__n12137), .Y(register__n12121) );
  INVx1_ASAP7_75t_R register___U7095 ( .A(register__net126178), .Y(register__net143255) );
  BUFx6f_ASAP7_75t_R register___U7096 ( .A(register__net63352), .Y(register__net126178) );
  INVx3_ASAP7_75t_R register___U7097 ( .A(register__n72), .Y(register__net62844) );
  BUFx4f_ASAP7_75t_R register___U7098 ( .A(register__n3645), .Y(register__n3469) );
  BUFx3_ASAP7_75t_R register___U7099 ( .A(register__n3645), .Y(register__n3470) );
  BUFx12f_ASAP7_75t_R register___U7100 ( .A(register__n1774), .Y(register__n3473) );
  BUFx12f_ASAP7_75t_R register___U7101 ( .A(register__n11904), .Y(register__n3480) );
  INVx6_ASAP7_75t_R register___U7102 ( .A(register__n3843), .Y(register__n6679) );
  INVx2_ASAP7_75t_R register___U7103 ( .A(register__n3481), .Y(register__n12428) );
  BUFx2_ASAP7_75t_R register___U7104 ( .A(register__n3485), .Y(register__n3484) );
  BUFx2_ASAP7_75t_R register___U7105 ( .A(register__n12871), .Y(register__n3485) );
  BUFx2_ASAP7_75t_R register___U7106 ( .A(register__n3487), .Y(register__n3486) );
  BUFx2_ASAP7_75t_R register___U7107 ( .A(register__n12985), .Y(register__n3487) );
  BUFx2_ASAP7_75t_R register___U7108 ( .A(register__n3489), .Y(register__n3488) );
  BUFx2_ASAP7_75t_R register___U7109 ( .A(register__n13220), .Y(register__n3489) );
  BUFx2_ASAP7_75t_R register___U7110 ( .A(register__n3491), .Y(register__n3490) );
  BUFx2_ASAP7_75t_R register___U7111 ( .A(register__n13010), .Y(register__n3491) );
  BUFx2_ASAP7_75t_R register___U7112 ( .A(register__n7070), .Y(register__n3494) );
  BUFx3_ASAP7_75t_R register___U7113 ( .A(register__n3496), .Y(register__n3495) );
  BUFx2_ASAP7_75t_R register___U7114 ( .A(register__n10559), .Y(register__n3496) );
  BUFx12f_ASAP7_75t_R register___U7115 ( .A(register__n6265), .Y(register__n12067) );
  INVx2_ASAP7_75t_R register___U7116 ( .A(register__net102926), .Y(register__net142928) );
  BUFx12f_ASAP7_75t_R register___U7117 ( .A(register__net145245), .Y(register__net102926) );
  BUFx3_ASAP7_75t_R register___U7118 ( .A(register__n8458), .Y(register__n3499) );
  BUFx6f_ASAP7_75t_R register___U7119 ( .A(register__n8457), .Y(register__n9296) );
  BUFx4f_ASAP7_75t_R register___U7120 ( .A(register__n3499), .Y(register__n8457) );
  BUFx6f_ASAP7_75t_R register___U7121 ( .A(register__n12040), .Y(register__n12025) );
  BUFx4f_ASAP7_75t_R register___U7122 ( .A(register__n4866), .Y(register__n12040) );
  INVx2_ASAP7_75t_R register___U7123 ( .A(register__n12380), .Y(register__n12366) );
  BUFx4f_ASAP7_75t_R register___U7124 ( .A(register__n3299), .Y(register__n12380) );
  OA22x2_ASAP7_75t_R register___U7125 ( .A1(register__n12150), .A2(register__n1974), .B1(register__n10132), .B2(register__n2829), 
        .Y(register__n12905) );
  INVx6_ASAP7_75t_R register___U7126 ( .A(register__n12161), .Y(register__n12150) );
  INVx4_ASAP7_75t_R register___U7127 ( .A(register__n12216), .Y(register__n12200) );
  BUFx12f_ASAP7_75t_R register___U7128 ( .A(register__n7257), .Y(register__n12096) );
  BUFx12f_ASAP7_75t_R register___U7129 ( .A(register__net141443), .Y(register__net142813) );
  BUFx12f_ASAP7_75t_R register___U7130 ( .A(register__net121464), .Y(register__net142807) );
  BUFx12f_ASAP7_75t_R register___U7131 ( .A(register__n3676), .Y(register__n3505) );
  BUFx12f_ASAP7_75t_R register___U7132 ( .A(register__n3676), .Y(register__n3506) );
  INVx5_ASAP7_75t_R register___U7133 ( .A(register__net64974), .Y(register__net64944) );
  INVx6_ASAP7_75t_R register___U7134 ( .A(register__net63208), .Y(register__net63174) );
  INVx6_ASAP7_75t_R register___U7135 ( .A(register__net138884), .Y(register__net63348) );
  INVx6_ASAP7_75t_R register___U7136 ( .A(register__n12074), .Y(register__n12063) );
  BUFx2_ASAP7_75t_R register___U7137 ( .A(register__n3519), .Y(register__n3518) );
  BUFx2_ASAP7_75t_R register___U7138 ( .A(register__n12995), .Y(register__n3519) );
  BUFx2_ASAP7_75t_R register___U7139 ( .A(register__n3521), .Y(register__n3520) );
  BUFx3_ASAP7_75t_R register___U7140 ( .A(register__n3523), .Y(register__n3522) );
  BUFx2_ASAP7_75t_R register___U7141 ( .A(register__n10809), .Y(register__n3523) );
  BUFx3_ASAP7_75t_R register___U7142 ( .A(register__n3526), .Y(register__n3525) );
  BUFx2_ASAP7_75t_R register___U7143 ( .A(register__n10808), .Y(register__n3526) );
  BUFx3_ASAP7_75t_R register___U7144 ( .A(register__n3528), .Y(register__n3527) );
  BUFx2_ASAP7_75t_R register___U7145 ( .A(register__n10745), .Y(register__n3528) );
  BUFx3_ASAP7_75t_R register___U7146 ( .A(register__n10746), .Y(register__n3529) );
  BUFx2_ASAP7_75t_R register___U7147 ( .A(register__n4977), .Y(register__n3530) );
  BUFx12f_ASAP7_75t_R register___U7148 ( .A(register__n3532), .Y(register__n3531) );
  BUFx6f_ASAP7_75t_R register___U7149 ( .A(register__n4577), .Y(register__n3533) );
  INVx3_ASAP7_75t_R register___U7150 ( .A(register__net62878), .Y(register__net62842) );
  BUFx2_ASAP7_75t_R register___U7151 ( .A(register__net64760), .Y(register__net142376) );
  INVx2_ASAP7_75t_R register___U7152 ( .A(register__net64792), .Y(register__net64760) );
  BUFx12f_ASAP7_75t_R register___U7153 ( .A(register__net137456), .Y(register__net142360) );
  BUFx12f_ASAP7_75t_R register___U7154 ( .A(register__n4771), .Y(register__n3538) );
  BUFx12f_ASAP7_75t_R register___U7155 ( .A(register__n3514), .Y(register__n3542) );
  BUFx12f_ASAP7_75t_R register___U7156 ( .A(register__n4198), .Y(register__n3544) );
  BUFx12f_ASAP7_75t_R register___U7157 ( .A(register__n3515), .Y(register__n3545) );
  BUFx2_ASAP7_75t_R register___U7158 ( .A(register__n3553), .Y(register__n3552) );
  BUFx2_ASAP7_75t_R register___U7159 ( .A(register__n12593), .Y(register__n3553) );
  BUFx2_ASAP7_75t_R register___U7160 ( .A(register__n3557), .Y(register__n3556) );
  BUFx2_ASAP7_75t_R register___U7161 ( .A(register__n12987), .Y(register__n3557) );
  BUFx2_ASAP7_75t_R register___U7162 ( .A(register__n3559), .Y(register__n3558) );
  OA22x2_ASAP7_75t_R register___U7163 ( .A1(register__net64336), .A2(register__n1755), .B1(register__net90673), .B2(
        n3334), .Y(register__n13136) );
  OA22x2_ASAP7_75t_R register___U7164 ( .A1(register__n11956), .A2(register__n3343), .B1(register__n9296), .B2(register__n11878), 
        .Y(register__n12978) );
  INVx1_ASAP7_75t_R register___U7165 ( .A(register__n3051), .Y(register__n3563) );
  INVx3_ASAP7_75t_R register___U7166 ( .A(register__n12274), .Y(register__n12260) );
  BUFx12f_ASAP7_75t_R register___U7167 ( .A(register__n3420), .Y(register__n4836) );
  BUFx12f_ASAP7_75t_R register___U7168 ( .A(register__n3679), .Y(register__n3565) );
  BUFx12f_ASAP7_75t_R register___U7169 ( .A(register__net140614), .Y(register__net141991) );
  BUFx12f_ASAP7_75t_R register___U7170 ( .A(register__net140260), .Y(register__net141985) );
  BUFx12f_ASAP7_75t_R register___U7171 ( .A(register__n3567), .Y(register__n3566) );
  BUFx12f_ASAP7_75t_R register___U7172 ( .A(register__n4474), .Y(register__n3567) );
  BUFx12f_ASAP7_75t_R register___U7173 ( .A(register__n3726), .Y(register__n3570) );
  BUFx12f_ASAP7_75t_R register___U7174 ( .A(register__net140272), .Y(register__net141957) );
  BUFx12f_ASAP7_75t_R register___U7175 ( .A(register__n11758), .Y(register__n3572) );
  INVx6_ASAP7_75t_R register___U7176 ( .A(register__n3595), .Y(register__n11926) );
  BUFx2_ASAP7_75t_R register___U7177 ( .A(register__n3574), .Y(register__n3573) );
  BUFx2_ASAP7_75t_R register___U7178 ( .A(register__n12725), .Y(register__n3574) );
  BUFx2_ASAP7_75t_R register___U7179 ( .A(register__n3576), .Y(register__n3575) );
  BUFx2_ASAP7_75t_R register___U7180 ( .A(register__n12743), .Y(register__n3576) );
  BUFx2_ASAP7_75t_R register___U7181 ( .A(register__n3578), .Y(register__n3577) );
  BUFx2_ASAP7_75t_R register___U7182 ( .A(register__n3580), .Y(register__n3579) );
  BUFx2_ASAP7_75t_R register___U7183 ( .A(register__n3584), .Y(register__n3583) );
  BUFx2_ASAP7_75t_R register___U7184 ( .A(register__n12872), .Y(register__n3584) );
  BUFx2_ASAP7_75t_R register___U7185 ( .A(register__n3586), .Y(register__n3585) );
  BUFx2_ASAP7_75t_R register___U7186 ( .A(register__n13012), .Y(register__n3586) );
  INVx4_ASAP7_75t_R register___U7187 ( .A(register__n3322), .Y(register__n12290) );
  BUFx2_ASAP7_75t_R register___U7188 ( .A(register__n3588), .Y(register__n3587) );
  BUFx2_ASAP7_75t_R register___U7189 ( .A(register__n3590), .Y(register__n3589) );
  OA22x2_ASAP7_75t_R register___U7190 ( .A1(register__net64672), .A2(register__n1266), .B1(register__n9762), .B2(register__n3334), 
        .Y(register__n13140) );
  OA22x2_ASAP7_75t_R register___U7191 ( .A1(register__net64684), .A2(register__n100), .B1(register__n9297), .B2(register__n11772), 
        .Y(register__n12972) );
  INVx4_ASAP7_75t_R register___U7192 ( .A(register__n12413), .Y(register__n12402) );
  BUFx3_ASAP7_75t_R register___U7193 ( .A(register__net62850), .Y(register__net141519) );
  BUFx12f_ASAP7_75t_R register___U7194 ( .A(register__n3598), .Y(register__n3596) );
  BUFx12f_ASAP7_75t_R register___U7195 ( .A(register__n3453), .Y(register__n3597) );
  BUFx12f_ASAP7_75t_R register___U7196 ( .A(register__n3878), .Y(register__n3598) );
  BUFx12f_ASAP7_75t_R register___U7197 ( .A(register__n12188), .Y(register__n3600) );
  BUFx12f_ASAP7_75t_R register___U7198 ( .A(register__net141491), .Y(register__net141489) );
  BUFx12f_ASAP7_75t_R register___U7199 ( .A(register__net64708), .Y(register__net141491) );
  BUFx12f_ASAP7_75t_R register___U7200 ( .A(register__net140266), .Y(register__net141466) );
  BUFx12f_ASAP7_75t_R register___U7201 ( .A(register__net144154), .Y(register__net62712) );
  BUFx12f_ASAP7_75t_R register___U7202 ( .A(register__n11809), .Y(register__n3605) );
  BUFx12f_ASAP7_75t_R register___U7203 ( .A(register__net102924), .Y(register__net141443) );
  BUFx12f_ASAP7_75t_R register___U7204 ( .A(register__net142813), .Y(register__net64888) );
  BUFx12f_ASAP7_75t_R register___U7205 ( .A(register__n11866), .Y(register__n3606) );
  INVx6_ASAP7_75t_R register___U7206 ( .A(register__net136862), .Y(register__net62828) );
  INVx6_ASAP7_75t_R register___U7207 ( .A(register__net136861), .Y(register__net62830) );
  BUFx12f_ASAP7_75t_R register___U7208 ( .A(register__net139024), .Y(register__net63016) );
  BUFx2_ASAP7_75t_R register___U7209 ( .A(register__n3608), .Y(register__n3607) );
  BUFx2_ASAP7_75t_R register___U7210 ( .A(register__n3614), .Y(register__n3613) );
  BUFx2_ASAP7_75t_R register___U7211 ( .A(register__n12874), .Y(register__n3614) );
  BUFx2_ASAP7_75t_R register___U7212 ( .A(register__n3616), .Y(register__n3615) );
  BUFx3_ASAP7_75t_R register___U7213 ( .A(register__n3618), .Y(register__n3617) );
  BUFx2_ASAP7_75t_R register___U7214 ( .A(register__n11045), .Y(register__n3618) );
  BUFx3_ASAP7_75t_R register___U7215 ( .A(register__n3620), .Y(register__n3619) );
  BUFx2_ASAP7_75t_R register___U7216 ( .A(register__n10579), .Y(register__n3620) );
  BUFx3_ASAP7_75t_R register___U7217 ( .A(register__n10576), .Y(register__n3621) );
  BUFx3_ASAP7_75t_R register___U7218 ( .A(register__n3623), .Y(register__n3622) );
  BUFx2_ASAP7_75t_R register___U7219 ( .A(register__n10578), .Y(register__n3623) );
  BUFx3_ASAP7_75t_R register___U7220 ( .A(register__n3625), .Y(register__n3624) );
  BUFx2_ASAP7_75t_R register___U7221 ( .A(register__n11109), .Y(register__n3625) );
  BUFx3_ASAP7_75t_R register___U7222 ( .A(register__n3627), .Y(register__n3626) );
  BUFx2_ASAP7_75t_R register___U7223 ( .A(register__n11111), .Y(register__n3627) );
  BUFx12f_ASAP7_75t_R register___U7224 ( .A(register__n12127), .Y(register__n3629) );
  INVx6_ASAP7_75t_R register___U7225 ( .A(register__net63210), .Y(register__net63180) );
  BUFx3_ASAP7_75t_R register___U7226 ( .A(register__n3631), .Y(register__n3630) );
  BUFx2_ASAP7_75t_R register___U7227 ( .A(register__n10793), .Y(register__n3631) );
  BUFx3_ASAP7_75t_R register___U7228 ( .A(register__n3636), .Y(register__n3635) );
  BUFx2_ASAP7_75t_R register___U7229 ( .A(register__n10790), .Y(register__n3636) );
  BUFx3_ASAP7_75t_R register___U7230 ( .A(register__n3638), .Y(register__n3637) );
  BUFx2_ASAP7_75t_R register___U7231 ( .A(Reg_data[661]), .Y(register__n3638) );
  BUFx3_ASAP7_75t_R register___U7232 ( .A(register__net141143), .Y(register__net141142) );
  BUFx2_ASAP7_75t_R register___U7233 ( .A(Reg_data[459]), .Y(register__net141143) );
  OA22x2_ASAP7_75t_R register___U7234 ( .A1(register__net63166), .A2(register__n100), .B1(register__net110124), .B2(
        n3301), .Y(register__n12954) );
  INVx1_ASAP7_75t_R register___U7235 ( .A(register__n3045), .Y(register__n3639) );
  OA22x2_ASAP7_75t_R register___U7236 ( .A1(register__net64420), .A2(register__n1755), .B1(register__net103467), .B2(
        n3821), .Y(register__n13137) );
  INVx1_ASAP7_75t_R register___U7237 ( .A(register__n3197), .Y(register__n3640) );
  INVx1_ASAP7_75t_R register___U7238 ( .A(register__n3040), .Y(register__n3642) );
  INVx1_ASAP7_75t_R register___U7239 ( .A(register__n10767), .Y(register__n3643) );
  BUFx4f_ASAP7_75t_R register___U7240 ( .A(register__n11992), .Y(register__n3644) );
  INVx3_ASAP7_75t_R register___U7241 ( .A(register__n12414), .Y(register__n12403) );
  BUFx12f_ASAP7_75t_R register___U7242 ( .A(register__n4197), .Y(register__n3646) );
  BUFx12f_ASAP7_75t_R register___U7243 ( .A(register__n12265), .Y(register__n3648) );
  BUFx12f_ASAP7_75t_R register___U7244 ( .A(register__n3731), .Y(register__n3649) );
  BUFx12f_ASAP7_75t_R register___U7245 ( .A(register__net143489), .Y(register__net141040) );
  BUFx12f_ASAP7_75t_R register___U7246 ( .A(register__net64476), .Y(register__net141026) );
  BUFx12f_ASAP7_75t_R register___U7247 ( .A(register__n12163), .Y(register__n3650) );
  BUFx4f_ASAP7_75t_R register___U7248 ( .A(register__n6680), .Y(register__n12134) );
  BUFx2_ASAP7_75t_R register___U7249 ( .A(register__n3654), .Y(register__n3653) );
  BUFx2_ASAP7_75t_R register___U7250 ( .A(register__n12642), .Y(register__n3654) );
  BUFx2_ASAP7_75t_R register___U7251 ( .A(register__n3658), .Y(register__n3657) );
  BUFx2_ASAP7_75t_R register___U7252 ( .A(register__n12820), .Y(register__n3658) );
  BUFx2_ASAP7_75t_R register___U7253 ( .A(register__n3662), .Y(register__n3661) );
  OA22x2_ASAP7_75t_R register___U7254 ( .A1(register__n12370), .A2(register__n3343), .B1(register__n6896), .B2(register__n3278), 
        .Y(register__n12957) );
  INVx1_ASAP7_75t_R register___U7255 ( .A(register__n2830), .Y(register__n3664) );
  BUFx6f_ASAP7_75t_R register___U7256 ( .A(register__n12003), .Y(register__n11987) );
  BUFx12f_ASAP7_75t_R register___U7257 ( .A(register__net91738), .Y(register__net140686) );
  INVx2_ASAP7_75t_R register___U7258 ( .A(register__n12413), .Y(register__n12397) );
  BUFx12f_ASAP7_75t_R register___U7259 ( .A(register__net64060), .Y(register__net140674) );
  BUFx12f_ASAP7_75t_R register___U7260 ( .A(register__net140665), .Y(register__net140663) );
  BUFx12f_ASAP7_75t_R register___U7261 ( .A(register__n11936), .Y(register__n3670) );
  BUFx12f_ASAP7_75t_R register___U7262 ( .A(register__n3703), .Y(register__n3671) );
  BUFx12f_ASAP7_75t_R register___U7263 ( .A(register__n3703), .Y(register__n3672) );
  BUFx12f_ASAP7_75t_R register___U7264 ( .A(register__n5502), .Y(register__n3674) );
  BUFx12f_ASAP7_75t_R register___U7265 ( .A(register__n11836), .Y(register__n3676) );
  BUFx4f_ASAP7_75t_R register___U7266 ( .A(register__n12182), .Y(register__n3677) );
  BUFx12f_ASAP7_75t_R register___U7267 ( .A(register__n12182), .Y(register__n3678) );
  BUFx12f_ASAP7_75t_R register___U7268 ( .A(register__net64782), .Y(register__net140614) );
  BUFx12f_ASAP7_75t_R register___U7269 ( .A(register__n12078), .Y(register__n3679) );
  BUFx12f_ASAP7_75t_R register___U7270 ( .A(register__net100797), .Y(register__net140597) );
  BUFx12f_ASAP7_75t_R register___U7271 ( .A(register__net143516), .Y(register__net62704) );
  INVx6_ASAP7_75t_R register___U7272 ( .A(register__n3728), .Y(register__n12458) );
  BUFx2_ASAP7_75t_R register___U7273 ( .A(register__n3683), .Y(register__n3682) );
  BUFx2_ASAP7_75t_R register___U7274 ( .A(register__n12643), .Y(register__n3683) );
  BUFx2_ASAP7_75t_R register___U7275 ( .A(register__n3685), .Y(register__n3684) );
  BUFx3_ASAP7_75t_R register___U7276 ( .A(register__net140428), .Y(register__net140427) );
  BUFx2_ASAP7_75t_R register___U7277 ( .A(Reg_data[293]), .Y(register__net140428) );
  BUFx3_ASAP7_75t_R register___U7278 ( .A(register__n3692), .Y(register__n3691) );
  BUFx2_ASAP7_75t_R register___U7279 ( .A(Reg_data[291]), .Y(register__n3692) );
  BUFx3_ASAP7_75t_R register___U7280 ( .A(register__n3694), .Y(register__n3693) );
  BUFx2_ASAP7_75t_R register___U7281 ( .A(Reg_data[289]), .Y(register__n3694) );
  BUFx3_ASAP7_75t_R register___U7282 ( .A(register__net140416), .Y(register__net140415) );
  BUFx2_ASAP7_75t_R register___U7283 ( .A(Reg_data[312]), .Y(register__net140416) );
  BUFx3_ASAP7_75t_R register___U7284 ( .A(register__n3696), .Y(register__n3695) );
  BUFx2_ASAP7_75t_R register___U7285 ( .A(Reg_data[297]), .Y(register__n3696) );
  BUFx3_ASAP7_75t_R register___U7286 ( .A(register__n3698), .Y(register__n3697) );
  BUFx2_ASAP7_75t_R register___U7287 ( .A(Reg_data[315]), .Y(register__n3698) );
  OA22x2_ASAP7_75t_R register___U7288 ( .A1(register__net64342), .A2(register__n100), .B1(register__net110088), .B2(
        n11771), .Y(register__n12968) );
  BUFx4f_ASAP7_75t_R register___U7289 ( .A(register__n11986), .Y(register__n3700) );
  INVx3_ASAP7_75t_R register___U7290 ( .A(register__n12207), .Y(register__n12192) );
  BUFx12f_ASAP7_75t_R register___U7291 ( .A(register__net102923), .Y(register__net64882) );
  BUFx12f_ASAP7_75t_R register___U7292 ( .A(register__n3844), .Y(register__n3703) );
  BUFx12f_ASAP7_75t_R register___U7293 ( .A(register__net139862), .Y(register__net140298) );
  BUFx12f_ASAP7_75t_R register___U7294 ( .A(register__n12243), .Y(register__n3705) );
  BUFx12f_ASAP7_75t_R register___U7295 ( .A(register__net140639), .Y(register__net140283) );
  BUFx12f_ASAP7_75t_R register___U7296 ( .A(register__net140640), .Y(register__net140284) );
  BUFx12f_ASAP7_75t_R register___U7297 ( .A(register__n3707), .Y(register__n3706) );
  BUFx12f_ASAP7_75t_R register___U7298 ( .A(register__n5171), .Y(register__n3707) );
  BUFx12f_ASAP7_75t_R register___U7299 ( .A(register__net141956), .Y(register__net140271) );
  BUFx12f_ASAP7_75t_R register___U7300 ( .A(register__net125383), .Y(register__net140272) );
  BUFx12f_ASAP7_75t_R register___U7301 ( .A(register__net63372), .Y(register__net140266) );
  BUFx12f_ASAP7_75t_R register___U7302 ( .A(register__net129617), .Y(register__net140260) );
  BUFx2_ASAP7_75t_R register___U7303 ( .A(register__n3713), .Y(register__n3712) );
  BUFx2_ASAP7_75t_R register___U7304 ( .A(register__n12645), .Y(register__n3713) );
  AND4x1_ASAP7_75t_R register___U7305 ( .A(register__n10611), .B(register__n10612), .C(register__n866), .D(register__n10613), .Y(
        n8586) );
  OA22x2_ASAP7_75t_R register___U7306 ( .A1(register__n12051), .A2(register__n100), .B1(register__n6619), .B2(register__n1918), 
        .Y(register__n12971) );
  OA22x2_ASAP7_75t_R register___U7307 ( .A1(register__net64416), .A2(register__n11868), .B1(register__net101049), .B2(
        n3275), .Y(register__n13277) );
  OA22x2_ASAP7_75t_R register___U7308 ( .A1(register__net63168), .A2(register__n1973), .B1(register__net90017), .B2(
        n11798), .Y(register__n12894) );
  BUFx6f_ASAP7_75t_R register___U7309 ( .A(register__n12001), .Y(register__n11984) );
  INVx3_ASAP7_75t_R register___U7310 ( .A(register__n11984), .Y(register__n3723) );
  BUFx4f_ASAP7_75t_R register___U7311 ( .A(register__n12219), .Y(register__n3724) );
  BUFx12f_ASAP7_75t_R register___U7312 ( .A(register__n12219), .Y(register__n3725) );
  INVx2_ASAP7_75t_R register___U7313 ( .A(register__n3725), .Y(register__n5684) );
  INVx4_ASAP7_75t_R register___U7314 ( .A(register__net63044), .Y(register__net63008) );
  BUFx12f_ASAP7_75t_R register___U7315 ( .A(register__net144561), .Y(register__net63044) );
  BUFx12f_ASAP7_75t_R register___U7316 ( .A(register__n3504), .Y(register__n11978) );
  BUFx12f_ASAP7_75t_R register___U7317 ( .A(register__n5353), .Y(register__n3728) );
  BUFx12f_ASAP7_75t_R register___U7318 ( .A(register__net141048), .Y(register__net139892) );
  BUFx12f_ASAP7_75t_R register___U7319 ( .A(register__n3649), .Y(register__n3729) );
  BUFx12f_ASAP7_75t_R register___U7320 ( .A(register__n3649), .Y(register__n3730) );
  BUFx12f_ASAP7_75t_R register___U7321 ( .A(register__n12442), .Y(register__n3731) );
  BUFx12f_ASAP7_75t_R register___U7322 ( .A(register__net64034), .Y(register__net64046) );
  BUFx12f_ASAP7_75t_R register___U7323 ( .A(register__net140298), .Y(register__net139860) );
  BUFx12f_ASAP7_75t_R register___U7324 ( .A(register__net64702), .Y(register__net139862) );
  BUFx12f_ASAP7_75t_R register___U7325 ( .A(register__n12247), .Y(register__n3733) );
  INVx6_ASAP7_75t_R register___U7326 ( .A(register__n12359), .Y(register__n12341) );
  BUFx12f_ASAP7_75t_R register___U7327 ( .A(register__n3565), .Y(register__n12076) );
  BUFx2_ASAP7_75t_R register___U7328 ( .A(register__net35927), .Y(register__net139812) );
  BUFx2_ASAP7_75t_R register___U7329 ( .A(register__n3739), .Y(register__n3738) );
  BUFx2_ASAP7_75t_R register___U7330 ( .A(register__n3745), .Y(register__n3744) );
  BUFx2_ASAP7_75t_R register___U7331 ( .A(register__n12644), .Y(register__n3745) );
  BUFx3_ASAP7_75t_R register___U7332 ( .A(register__n3748), .Y(register__n3747) );
  BUFx2_ASAP7_75t_R register___U7333 ( .A(Reg_data[305]), .Y(register__n3748) );
  BUFx3_ASAP7_75t_R register___U7334 ( .A(register__n3750), .Y(register__n3749) );
  BUFx2_ASAP7_75t_R register___U7335 ( .A(Reg_data[307]), .Y(register__n3750) );
  OA22x2_ASAP7_75t_R register___U7336 ( .A1(register__n11927), .A2(register__n3343), .B1(register__n6909), .B2(register__n11880), 
        .Y(register__n12979) );
  OA22x2_ASAP7_75t_R register___U7337 ( .A1(register__n12112), .A2(register__n1408), .B1(register__n8155), .B2(register__n2882), 
        .Y(register__n13276) );
  OA22x2_ASAP7_75t_R register___U7338 ( .A1(register__n12118), .A2(register__n1973), .B1(register__n10157), .B2(register__n11882), 
        .Y(register__n12906) );
  INVx1_ASAP7_75t_R register___U7339 ( .A(register__n3006), .Y(register__n3753) );
  BUFx12f_ASAP7_75t_R register___U7340 ( .A(register__n4842), .Y(register__n11903) );
  BUFx12f_ASAP7_75t_R register___U7341 ( .A(register__n3568), .Y(register__n4728) );
  BUFx12f_ASAP7_75t_R register___U7342 ( .A(register__net141040), .Y(register__net64974) );
  BUFx12f_ASAP7_75t_R register___U7343 ( .A(register__net141039), .Y(register__net64966) );
  BUFx2_ASAP7_75t_R register___U7344 ( .A(register__n3758), .Y(register__n3757) );
  BUFx2_ASAP7_75t_R register___U7345 ( .A(register__n12537), .Y(register__n3758) );
  BUFx2_ASAP7_75t_R register___U7346 ( .A(register__n3761), .Y(register__n3760) );
  BUFx2_ASAP7_75t_R register___U7347 ( .A(register__n12544), .Y(register__n3761) );
  BUFx2_ASAP7_75t_R register___U7348 ( .A(register__n3763), .Y(register__n3762) );
  BUFx2_ASAP7_75t_R register___U7349 ( .A(register__n12744), .Y(register__n3763) );
  BUFx2_ASAP7_75t_R register___U7350 ( .A(register__n3766), .Y(register__n3765) );
  BUFx2_ASAP7_75t_R register___U7351 ( .A(register__n3768), .Y(register__n3767) );
  BUFx2_ASAP7_75t_R register___U7352 ( .A(register__n13093), .Y(register__n3768) );
  BUFx2_ASAP7_75t_R register___U7353 ( .A(register__n3774), .Y(register__n3773) );
  BUFx2_ASAP7_75t_R register___U7354 ( .A(register__n12817), .Y(register__n3774) );
  BUFx2_ASAP7_75t_R register___U7355 ( .A(register__n3776), .Y(register__n3775) );
  BUFx2_ASAP7_75t_R register___U7356 ( .A(register__n3778), .Y(register__n3777) );
  BUFx2_ASAP7_75t_R register___U7357 ( .A(register__n12821), .Y(register__n3778) );
  BUFx2_ASAP7_75t_R register___U7358 ( .A(register__n3780), .Y(register__n3779) );
  BUFx2_ASAP7_75t_R register___U7359 ( .A(register__n12724), .Y(register__n3785) );
  BUFx12f_ASAP7_75t_R register___U7360 ( .A(register__n3447), .Y(register__n12300) );
  BUFx4f_ASAP7_75t_R register___U7361 ( .A(register__n3791), .Y(register__n3790) );
  BUFx3_ASAP7_75t_R register___U7362 ( .A(register__n8379), .Y(register__n3791) );
  BUFx6f_ASAP7_75t_R register___U7363 ( .A(register__n3790), .Y(register__n10157) );
  BUFx3_ASAP7_75t_R register___U7364 ( .A(register__net139227), .Y(register__net139226) );
  BUFx2_ASAP7_75t_R register___U7365 ( .A(Reg_data[569]), .Y(register__net139227) );
  BUFx3_ASAP7_75t_R register___U7366 ( .A(register__n3795), .Y(register__n3794) );
  BUFx2_ASAP7_75t_R register___U7367 ( .A(Reg_data[565]), .Y(register__n3795) );
  BUFx3_ASAP7_75t_R register___U7368 ( .A(register__n3797), .Y(register__n3796) );
  BUFx2_ASAP7_75t_R register___U7369 ( .A(Reg_data[564]), .Y(register__n3797) );
  BUFx3_ASAP7_75t_R register___U7370 ( .A(register__n3799), .Y(register__n3798) );
  BUFx2_ASAP7_75t_R register___U7371 ( .A(Reg_data[562]), .Y(register__n3799) );
  BUFx3_ASAP7_75t_R register___U7372 ( .A(register__n3801), .Y(register__n3800) );
  BUFx2_ASAP7_75t_R register___U7373 ( .A(Reg_data[560]), .Y(register__n3801) );
  BUFx3_ASAP7_75t_R register___U7374 ( .A(register__net139207), .Y(register__net139206) );
  BUFx2_ASAP7_75t_R register___U7375 ( .A(Reg_data[550]), .Y(register__net139207) );
  BUFx3_ASAP7_75t_R register___U7376 ( .A(register__net139203), .Y(register__net139202) );
  BUFx2_ASAP7_75t_R register___U7377 ( .A(Reg_data[549]), .Y(register__net139203) );
  BUFx3_ASAP7_75t_R register___U7378 ( .A(register__n3803), .Y(register__n3802) );
  BUFx2_ASAP7_75t_R register___U7379 ( .A(Reg_data[546]), .Y(register__n3803) );
  BUFx3_ASAP7_75t_R register___U7380 ( .A(register__n3805), .Y(register__n3804) );
  BUFx2_ASAP7_75t_R register___U7381 ( .A(Reg_data[544]), .Y(register__n3805) );
  BUFx3_ASAP7_75t_R register___U7382 ( .A(register__n3807), .Y(register__n3806) );
  BUFx2_ASAP7_75t_R register___U7383 ( .A(Reg_data[553]), .Y(register__n3807) );
  BUFx3_ASAP7_75t_R register___U7384 ( .A(register__net139187), .Y(register__net139186) );
  BUFx2_ASAP7_75t_R register___U7385 ( .A(Reg_data[555]), .Y(register__net139187) );
  BUFx3_ASAP7_75t_R register___U7386 ( .A(register__net139183), .Y(register__net139182) );
  BUFx2_ASAP7_75t_R register___U7387 ( .A(Reg_data[568]), .Y(register__net139183) );
  BUFx3_ASAP7_75t_R register___U7388 ( .A(register__net139179), .Y(register__net139178) );
  BUFx2_ASAP7_75t_R register___U7389 ( .A(Reg_data[559]), .Y(register__net139179) );
  BUFx3_ASAP7_75t_R register___U7390 ( .A(register__n3809), .Y(register__n3808) );
  BUFx2_ASAP7_75t_R register___U7391 ( .A(Reg_data[551]), .Y(register__n3809) );
  BUFx3_ASAP7_75t_R register___U7392 ( .A(register__n3811), .Y(register__n3810) );
  BUFx2_ASAP7_75t_R register___U7393 ( .A(Reg_data[558]), .Y(register__n3811) );
  BUFx3_ASAP7_75t_R register___U7394 ( .A(register__net139167), .Y(register__net139166) );
  BUFx2_ASAP7_75t_R register___U7395 ( .A(Reg_data[554]), .Y(register__net139167) );
  BUFx3_ASAP7_75t_R register___U7396 ( .A(register__n3813), .Y(register__n3812) );
  BUFx2_ASAP7_75t_R register___U7397 ( .A(Reg_data[563]), .Y(register__n3813) );
  BUFx3_ASAP7_75t_R register___U7398 ( .A(register__n3815), .Y(register__n3814) );
  BUFx2_ASAP7_75t_R register___U7399 ( .A(Reg_data[567]), .Y(register__n3815) );
  BUFx3_ASAP7_75t_R register___U7400 ( .A(register__n3817), .Y(register__n3816) );
  BUFx2_ASAP7_75t_R register___U7401 ( .A(Reg_data[570]), .Y(register__n3817) );
  BUFx3_ASAP7_75t_R register___U7402 ( .A(register__n3819), .Y(register__n3818) );
  BUFx2_ASAP7_75t_R register___U7403 ( .A(Reg_data[561]), .Y(register__n3819) );
  OA22x2_ASAP7_75t_R register___U7404 ( .A1(register__n12343), .A2(register__n3343), .B1(register__n6914), .B2(register__n2966), 
        .Y(register__n12958) );
  OA22x2_ASAP7_75t_R register___U7405 ( .A1(register__net63324), .A2(register__n1409), .B1(register__n6646), .B2(register__n3274), 
        .Y(register__n13269) );
  INVx4_ASAP7_75t_R register___U7406 ( .A(register__n12041), .Y(register__n4045) );
  BUFx12f_ASAP7_75t_R register___U7407 ( .A(register__net143491), .Y(register__net139023) );
  BUFx12f_ASAP7_75t_R register___U7408 ( .A(register__net143492), .Y(register__net139024) );
  BUFx12f_ASAP7_75t_R register___U7409 ( .A(register__net139016), .Y(register__net64478) );
  BUFx12f_ASAP7_75t_R register___U7410 ( .A(register__n11761), .Y(register__n3822) );
  INVx6_ASAP7_75t_R register___U7411 ( .A(register__net133742), .Y(register__net64348) );
  BUFx2_ASAP7_75t_R register___U7412 ( .A(register__n3825), .Y(register__n3824) );
  BUFx2_ASAP7_75t_R register___U7413 ( .A(register__n3827), .Y(register__n3826) );
  BUFx12f_ASAP7_75t_R register___U7414 ( .A(register__net142763), .Y(register__net138884) );
  BUFx12f_ASAP7_75t_R register___U7415 ( .A(register__net142763), .Y(register__net138885) );
  BUFx12f_ASAP7_75t_R register___U7416 ( .A(register__n3503), .Y(register__n3833) );
  BUFx12f_ASAP7_75t_R register___U7417 ( .A(register__n3833), .Y(register__n11979) );
  OA22x2_ASAP7_75t_R register___U7418 ( .A1(register__n12286), .A2(register__n101), .B1(register__n6955), .B2(register__n2854), 
        .Y(register__n12960) );
  OA22x2_ASAP7_75t_R register___U7419 ( .A1(register__n12396), .A2(register__n2851), .B1(register__n6663), .B2(register__n11869), 
        .Y(register__n13266) );
  INVx1_ASAP7_75t_R register___U7420 ( .A(register__n13266), .Y(register__n3834) );
  OA22x2_ASAP7_75t_R register___U7421 ( .A1(register__n12169), .A2(register__n1755), .B1(register__n7808), .B2(register__n3821), 
        .Y(register__n13133) );
  INVx1_ASAP7_75t_R register___U7422 ( .A(register__n3162), .Y(register__n3836) );
  OA22x2_ASAP7_75t_R register___U7423 ( .A1(register__net63252), .A2(register__n1973), .B1(register__net88504), .B2(
        n11791), .Y(register__n12895) );
  BUFx12f_ASAP7_75t_R register___U7424 ( .A(register__net64056), .Y(register__net64034) );
  BUFx12f_ASAP7_75t_R register___U7425 ( .A(register__net138596), .Y(register__net130079) );
  BUFx12f_ASAP7_75t_R register___U7426 ( .A(register__net138028), .Y(register__net138596) );
  BUFx12f_ASAP7_75t_R register___U7427 ( .A(register__n3876), .Y(register__n3840) );
  BUFx12f_ASAP7_75t_R register___U7428 ( .A(register__net138032), .Y(register__net138559) );
  BUFx12f_ASAP7_75t_R register___U7429 ( .A(register__n3283), .Y(register__n12359) );
  BUFx12f_ASAP7_75t_R register___U7430 ( .A(register__n3536), .Y(register__n3841) );
  BUFx12f_ASAP7_75t_R register___U7431 ( .A(register__n3534), .Y(register__n11939) );
  BUFx12f_ASAP7_75t_R register___U7432 ( .A(register__n3672), .Y(register__n3843) );
  BUFx12f_ASAP7_75t_R register___U7433 ( .A(register__n3848), .Y(register__n3846) );
  BUFx12f_ASAP7_75t_R register___U7434 ( .A(register__n3848), .Y(register__n3847) );
  BUFx12f_ASAP7_75t_R register___U7435 ( .A(register__n12015), .Y(register__n3848) );
  BUFx12f_ASAP7_75t_R register___U7436 ( .A(register__n12016), .Y(register__n12015) );
  BUFx3_ASAP7_75t_R register___U7437 ( .A(register__n3850), .Y(register__n3849) );
  BUFx2_ASAP7_75t_R register___U7438 ( .A(register__n11488), .Y(register__n3850) );
  BUFx3_ASAP7_75t_R register___U7439 ( .A(register__n3852), .Y(register__n3851) );
  BUFx2_ASAP7_75t_R register___U7440 ( .A(register__n11209), .Y(register__n3852) );
  BUFx2_ASAP7_75t_R register___U7441 ( .A(register__n3856), .Y(register__n3855) );
  BUFx2_ASAP7_75t_R register___U7442 ( .A(register__n12698), .Y(register__n3856) );
  BUFx2_ASAP7_75t_R register___U7443 ( .A(register__n3860), .Y(register__n3859) );
  BUFx2_ASAP7_75t_R register___U7444 ( .A(register__n13049), .Y(register__n3860) );
  BUFx2_ASAP7_75t_R register___U7445 ( .A(register__n5533), .Y(register__n3863) );
  BUFx3_ASAP7_75t_R register___U7446 ( .A(register__n3865), .Y(register__n3864) );
  BUFx2_ASAP7_75t_R register___U7447 ( .A(register__n11005), .Y(register__n3865) );
  BUFx12f_ASAP7_75t_R register___U7448 ( .A(register__n7610), .Y(register__n11972) );
  OA22x2_ASAP7_75t_R register___U7449 ( .A1(register__net64426), .A2(register__n100), .B1(register__net112283), .B2(
        n2844), .Y(register__n12969) );
  OA22x2_ASAP7_75t_R register___U7450 ( .A1(register__net63240), .A2(register__n1408), .B1(register__net100894), .B2(
        n2855), .Y(register__n13268) );
  OA22x2_ASAP7_75t_R register___U7451 ( .A1(register__n12252), .A2(register__n1755), .B1(register__n9688), .B2(register__n3821), 
        .Y(register__n13129) );
  OA22x2_ASAP7_75t_R register___U7452 ( .A1(register__n12371), .A2(register__n1974), .B1(register__n9969), .B2(register__n11790), 
        .Y(register__n12897) );
  BUFx2_ASAP7_75t_R register___U7453 ( .A(register__n5983), .Y(register__n3874) );
  BUFx2_ASAP7_75t_R register___U7454 ( .A(register__n6395), .Y(register__n3875) );
  BUFx12f_ASAP7_75t_R register___U7455 ( .A(register__n12438), .Y(register__n3876) );
  BUFx12f_ASAP7_75t_R register___U7456 ( .A(register__net138559), .Y(register__net138031) );
  BUFx12f_ASAP7_75t_R register___U7457 ( .A(register__net64712), .Y(register__net138032) );
  INVx6_ASAP7_75t_R register___U7458 ( .A(register__net138031), .Y(register__net64668) );
  BUFx12f_ASAP7_75t_R register___U7459 ( .A(register__n12335), .Y(register__n3878) );
  BUFx12f_ASAP7_75t_R register___U7460 ( .A(register__n3187), .Y(register__n11981) );
  BUFx12f_ASAP7_75t_R register___U7461 ( .A(register__n11971), .Y(register__n11980) );
  BUFx3_ASAP7_75t_R register___U7462 ( .A(register__n3881), .Y(register__n3880) );
  BUFx2_ASAP7_75t_R register___U7463 ( .A(register__n11608), .Y(register__n3881) );
  BUFx2_ASAP7_75t_R register___U7464 ( .A(register__n3885), .Y(register__n3884) );
  BUFx2_ASAP7_75t_R register___U7465 ( .A(register__n3894), .Y(register__n3893) );
  BUFx2_ASAP7_75t_R register___U7466 ( .A(register__n3896), .Y(register__n3895) );
  BUFx2_ASAP7_75t_R register___U7467 ( .A(register__n13206), .Y(register__n3896) );
  BUFx2_ASAP7_75t_R register___U7468 ( .A(register__n3898), .Y(register__n3897) );
  BUFx2_ASAP7_75t_R register___U7469 ( .A(register__n3902), .Y(register__n3901) );
  BUFx2_ASAP7_75t_R register___U7470 ( .A(register__n12789), .Y(register__n3902) );
  BUFx2_ASAP7_75t_R register___U7471 ( .A(register__n3905), .Y(register__n3904) );
  BUFx2_ASAP7_75t_R register___U7472 ( .A(register__n13215), .Y(register__n3905) );
  BUFx2_ASAP7_75t_R register___U7473 ( .A(register__n13042), .Y(register__n3907) );
  BUFx12f_ASAP7_75t_R register___U7474 ( .A(register__net146267), .Y(register__net137769) );
  OA22x2_ASAP7_75t_R register___U7475 ( .A1(register__net63248), .A2(register__n952), .B1(register__net88416), .B2(register__n959), .Y(register__n13016) );
  OA22x2_ASAP7_75t_R register___U7476 ( .A1(register__n12230), .A2(register__n101), .B1(register__n6668), .B2(register__n11779), 
        .Y(register__n12962) );
  INVx1_ASAP7_75t_R register___U7477 ( .A(register__n2865), .Y(register__n3910) );
  INVx1_ASAP7_75t_R register___U7478 ( .A(register__n2911), .Y(register__n3911) );
  OA22x2_ASAP7_75t_R register___U7479 ( .A1(register__net63160), .A2(register__n1755), .B1(register__net90813), .B2(
        n3821), .Y(register__n13122) );
  BUFx2_ASAP7_75t_R register___U7480 ( .A(register__n8662), .Y(register__n3913) );
  INVx4_ASAP7_75t_R register___U7481 ( .A(register__n12440), .Y(register__n12424) );
  BUFx3_ASAP7_75t_R register___U7482 ( .A(register__n10845), .Y(register__n3914) );
  BUFx4f_ASAP7_75t_R register___U7483 ( .A(register__n3914), .Y(register__n6779) );
  BUFx12f_ASAP7_75t_R register___U7484 ( .A(register__net63216), .Y(register__net63214) );
  BUFx12f_ASAP7_75t_R register___U7485 ( .A(register__n3671), .Y(register__n3916) );
  BUFx12f_ASAP7_75t_R register___U7486 ( .A(register__net128109), .Y(register__net137463) );
  BUFx12f_ASAP7_75t_R register___U7487 ( .A(register__n3847), .Y(register__n12008) );
  BUFx12f_ASAP7_75t_R register___U7488 ( .A(register__net142360), .Y(register__net64728) );
  BUFx12f_ASAP7_75t_R register___U7489 ( .A(register__net137418), .Y(register__net137417) );
  BUFx12f_ASAP7_75t_R register___U7490 ( .A(register__net143520), .Y(register__net63384) );
  BUFx12f_ASAP7_75t_R register___U7491 ( .A(register__net63384), .Y(register__net63372) );
  BUFx3_ASAP7_75t_R register___U7492 ( .A(register__n3921), .Y(register__n3920) );
  BUFx2_ASAP7_75t_R register___U7493 ( .A(register__n11507), .Y(register__n3921) );
  INVx6_ASAP7_75t_R register___U7494 ( .A(register__n11974), .Y(register__n11958) );
  BUFx12f_ASAP7_75t_R register___U7495 ( .A(register__n3412), .Y(register__n11974) );
  BUFx2_ASAP7_75t_R register___U7496 ( .A(register__n3923), .Y(register__n3922) );
  BUFx2_ASAP7_75t_R register___U7497 ( .A(register__n3929), .Y(register__n3928) );
  BUFx2_ASAP7_75t_R register___U7498 ( .A(register__n13332), .Y(register__n3929) );
  BUFx2_ASAP7_75t_R register___U7499 ( .A(register__n12875), .Y(register__n3931) );
  BUFx2_ASAP7_75t_R register___U7500 ( .A(register__n3933), .Y(register__n3932) );
  BUFx12f_ASAP7_75t_R register___U7501 ( .A(register__n5498), .Y(register__n3936) );
  INVx1_ASAP7_75t_R register___U7502 ( .A(register__n2862), .Y(register__n3941) );
  OA22x2_ASAP7_75t_R register___U7503 ( .A1(register__n12171), .A2(register__n100), .B1(register__n6982), .B2(register__n11780), 
        .Y(register__n12965) );
  INVx1_ASAP7_75t_R register___U7504 ( .A(register__n2869), .Y(register__n3943) );
  INVx1_ASAP7_75t_R register___U7505 ( .A(register__n2919), .Y(register__n3945) );
  OA22x2_ASAP7_75t_R register___U7506 ( .A1(register__n12314), .A2(register__n1755), .B1(register__n9686), .B2(register__n3336), 
        .Y(register__n13127) );
  BUFx12f_ASAP7_75t_R register___U7507 ( .A(register__net121482), .Y(register__net136861) );
  BUFx12f_ASAP7_75t_R register___U7508 ( .A(register__net62860), .Y(register__net136862) );
  BUFx12f_ASAP7_75t_R register___U7509 ( .A(register__net140663), .Y(register__net121482) );
  BUFx12f_ASAP7_75t_R register___U7510 ( .A(register__net142364), .Y(register__net64976) );
  BUFx2_ASAP7_75t_R register___U7511 ( .A(register__n3950), .Y(register__n3949) );
  BUFx2_ASAP7_75t_R register___U7512 ( .A(register__n12943), .Y(register__n3950) );
  BUFx2_ASAP7_75t_R register___U7513 ( .A(register__n3952), .Y(register__n3951) );
  BUFx2_ASAP7_75t_R register___U7514 ( .A(register__n13384), .Y(register__n3952) );
  BUFx2_ASAP7_75t_R register___U7515 ( .A(register__n3954), .Y(register__n3953) );
  BUFx2_ASAP7_75t_R register___U7516 ( .A(register__n13376), .Y(register__n3954) );
  BUFx2_ASAP7_75t_R register___U7517 ( .A(register__n3957), .Y(register__n3956) );
  BUFx2_ASAP7_75t_R register___U7518 ( .A(register__n3959), .Y(register__n3958) );
  BUFx2_ASAP7_75t_R register___U7519 ( .A(register__n13375), .Y(register__n3959) );
  BUFx2_ASAP7_75t_R register___U7520 ( .A(register__n3969), .Y(register__n3968) );
  BUFx2_ASAP7_75t_R register___U7521 ( .A(register__n3972), .Y(register__n3971) );
  BUFx2_ASAP7_75t_R register___U7522 ( .A(register__n13361), .Y(register__n3972) );
  BUFx2_ASAP7_75t_R register___U7523 ( .A(register__n12930), .Y(register__n3973) );
  INVx6_ASAP7_75t_R register___U7524 ( .A(register__n12244), .Y(register__n12231) );
  BUFx2_ASAP7_75t_R register___U7525 ( .A(register__n3979), .Y(register__n3978) );
  BUFx2_ASAP7_75t_R register___U7526 ( .A(register__n13358), .Y(register__n3979) );
  BUFx3_ASAP7_75t_R register___U7527 ( .A(register__n3981), .Y(register__n3980) );
  BUFx2_ASAP7_75t_R register___U7528 ( .A(register__n11334), .Y(register__n3981) );
  BUFx3_ASAP7_75t_R register___U7529 ( .A(register__n3983), .Y(register__n3982) );
  BUFx2_ASAP7_75t_R register___U7530 ( .A(register__n11336), .Y(register__n3983) );
  BUFx2_ASAP7_75t_R register___U7531 ( .A(register__n6148), .Y(register__n3984) );
  BUFx3_ASAP7_75t_R register___U7532 ( .A(register__n3986), .Y(register__n3985) );
  BUFx2_ASAP7_75t_R register___U7533 ( .A(register__n10942), .Y(register__n3986) );
  BUFx2_ASAP7_75t_R register___U7534 ( .A(register__n10583), .Y(register__n3987) );
  BUFx2_ASAP7_75t_R register___U7535 ( .A(register__n5700), .Y(register__n3988) );
  BUFx3_ASAP7_75t_R register___U7536 ( .A(register__n3990), .Y(register__n3989) );
  BUFx2_ASAP7_75t_R register___U7537 ( .A(register__n10580), .Y(register__n3990) );
  BUFx6f_ASAP7_75t_R register___U7538 ( .A(register__n12048), .Y(register__n3992) );
  AND4x1_ASAP7_75t_R register___U7539 ( .A(register__n11195), .B(register__n11196), .C(register__n11197), .D(register__n231), .Y(
        n7612) );
  INVx1_ASAP7_75t_R register___U7540 ( .A(register__n3657), .Y(register__n3995) );
  OA22x2_ASAP7_75t_R register___U7541 ( .A1(register__n12198), .A2(register__n3343), .B1(register__n6893), .B2(register__n3185), 
        .Y(register__n12963) );
  OA22x2_ASAP7_75t_R register___U7542 ( .A1(register__net63334), .A2(register__n956), .B1(register__n9764), .B2(register__n958), 
        .Y(register__n13017) );
  OA22x2_ASAP7_75t_R register___U7543 ( .A1(register__n12256), .A2(register__n1973), .B1(register__n9973), .B2(register__n11788), 
        .Y(register__n12901) );
  INVx1_ASAP7_75t_R register___U7544 ( .A(register__n2925), .Y(register__n3998) );
  BUFx12f_ASAP7_75t_R register___U7545 ( .A(register__net64710), .Y(register__net136275) );
  BUFx12f_ASAP7_75t_R register___U7546 ( .A(register__net127693), .Y(register__net136246) );
  BUFx3_ASAP7_75t_R register___U7547 ( .A(register__net127692), .Y(register__net136247) );
  BUFx4f_ASAP7_75t_R register___U7548 ( .A(register__net127693), .Y(register__net136248) );
  BUFx12f_ASAP7_75t_R register___U7549 ( .A(register__net136246), .Y(register__net64796) );
  OR2x2_ASAP7_75t_R register___U7550 ( .A(register__n5769), .B(register__n4002), .Y(register__n13203) );
  BUFx12f_ASAP7_75t_R register___U7551 ( .A(register__n3916), .Y(register__n12305) );
  BUFx2_ASAP7_75t_R register___U7552 ( .A(register__n5744), .Y(register__n4003) );
  BUFx12f_ASAP7_75t_R register___U7553 ( .A(register__net145051), .Y(register__net136187) );
  BUFx2_ASAP7_75t_R register___U7554 ( .A(register__n4006), .Y(register__n4005) );
  BUFx2_ASAP7_75t_R register___U7555 ( .A(register__n4010), .Y(register__n4009) );
  BUFx2_ASAP7_75t_R register___U7556 ( .A(register__n13197), .Y(register__n4010) );
  BUFx2_ASAP7_75t_R register___U7557 ( .A(register__n4012), .Y(register__n4011) );
  BUFx3_ASAP7_75t_R register___U7558 ( .A(register__n11487), .Y(register__n4015) );
  BUFx2_ASAP7_75t_R register___U7559 ( .A(register__n6407), .Y(register__n4018) );
  BUFx3_ASAP7_75t_R register___U7560 ( .A(register__n4020), .Y(register__n4019) );
  BUFx2_ASAP7_75t_R register___U7561 ( .A(register__n11486), .Y(register__n4020) );
  BUFx2_ASAP7_75t_R register___U7562 ( .A(register__n1071), .Y(register__n4021) );
  BUFx3_ASAP7_75t_R register___U7563 ( .A(register__n11114), .Y(register__n4025) );
  BUFx2_ASAP7_75t_R register___U7564 ( .A(register__n5928), .Y(register__n4026) );
  BUFx3_ASAP7_75t_R register___U7565 ( .A(register__n4028), .Y(register__n4027) );
  BUFx12f_ASAP7_75t_R register___U7566 ( .A(register__net74029), .Y(register__net74027) );
  INVx1_ASAP7_75t_R register___U7567 ( .A(register__n2898), .Y(register__n4038) );
  BUFx3_ASAP7_75t_R register___U7568 ( .A(register__net135779), .Y(register__net135778) );
  BUFx2_ASAP7_75t_R register___U7569 ( .A(Reg_data[153]), .Y(register__net135779) );
  BUFx3_ASAP7_75t_R register___U7570 ( .A(register__net135775), .Y(register__net135774) );
  BUFx2_ASAP7_75t_R register___U7571 ( .A(Reg_data[133]), .Y(register__net135775) );
  BUFx3_ASAP7_75t_R register___U7572 ( .A(register__n4040), .Y(register__n4039) );
  BUFx2_ASAP7_75t_R register___U7573 ( .A(Reg_data[132]), .Y(register__n4040) );
  BUFx3_ASAP7_75t_R register___U7574 ( .A(register__n4042), .Y(register__n4041) );
  BUFx2_ASAP7_75t_R register___U7575 ( .A(Reg_data[130]), .Y(register__n4042) );
  BUFx3_ASAP7_75t_R register___U7576 ( .A(register__net135763), .Y(register__net135762) );
  BUFx2_ASAP7_75t_R register___U7577 ( .A(Reg_data[143]), .Y(register__net135763) );
  BUFx3_ASAP7_75t_R register___U7578 ( .A(register__n4044), .Y(register__n4043) );
  BUFx2_ASAP7_75t_R register___U7579 ( .A(Reg_data[145]), .Y(register__n4044) );
  INVx2_ASAP7_75t_R register___U7580 ( .A(register__n12041), .Y(register__n12020) );
  OA22x2_ASAP7_75t_R register___U7581 ( .A1(register__n12142), .A2(register__n11730), .B1(register__n9523), .B2(register__n1164), 
        .Y(register__n13376) );
  INVx1_ASAP7_75t_R register___U7582 ( .A(register__n3953), .Y(register__n4046) );
  INVx6_ASAP7_75t_R register___U7583 ( .A(register__n12155), .Y(register__n12142) );
  OA22x2_ASAP7_75t_R register___U7584 ( .A1(register__n12151), .A2(register__n665), .B1(register__n8454), .B2(register__n81), .Y(
        n12818) );
  INVx1_ASAP7_75t_R register___U7585 ( .A(register__n3462), .Y(register__n4047) );
  INVx6_ASAP7_75t_R register___U7586 ( .A(register__net62696), .Y(register__net62652) );
  OA22x2_ASAP7_75t_R register___U7587 ( .A1(register__n12199), .A2(register__n1913), .B1(register__n8789), .B2(register__n11786), 
        .Y(register__n12903) );
  OA22x2_ASAP7_75t_R register___U7588 ( .A1(register__n12342), .A2(register__n952), .B1(register__n8807), .B2(register__n960), 
        .Y(register__n13019) );
  OA22x2_ASAP7_75t_R register___U7589 ( .A1(register__n12054), .A2(register__n1266), .B1(register__n7990), .B2(register__n3334), 
        .Y(register__n13139) );
  BUFx3_ASAP7_75t_R register___U7590 ( .A(register__n4051), .Y(register__n4050) );
  BUFx2_ASAP7_75t_R register___U7591 ( .A(register__n11250), .Y(register__n4051) );
  BUFx3_ASAP7_75t_R register___U7592 ( .A(register__n4053), .Y(register__n4052) );
  BUFx2_ASAP7_75t_R register___U7593 ( .A(register__n11396), .Y(register__n4053) );
  AO22x1_ASAP7_75t_R register___U7594 ( .A1(register__n9752), .A2(register__C6423_net61318), .B1(register__n8117), .B2(
        n1452), .Y(register__n11396) );
  INVx6_ASAP7_75t_R register___U7595 ( .A(register__n3733), .Y(register__n12236) );
  BUFx2_ASAP7_75t_R register___U7596 ( .A(register__n4055), .Y(register__n4054) );
  BUFx2_ASAP7_75t_R register___U7597 ( .A(register__n12873), .Y(register__n4055) );
  BUFx2_ASAP7_75t_R register___U7598 ( .A(register__n4057), .Y(register__n4056) );
  BUFx2_ASAP7_75t_R register___U7599 ( .A(register__n4059), .Y(register__n4058) );
  BUFx2_ASAP7_75t_R register___U7600 ( .A(register__n13262), .Y(register__n4059) );
  BUFx2_ASAP7_75t_R register___U7601 ( .A(register__n4063), .Y(register__n4062) );
  BUFx2_ASAP7_75t_R register___U7602 ( .A(register__n13329), .Y(register__n4063) );
  BUFx2_ASAP7_75t_R register___U7603 ( .A(register__n4065), .Y(register__n4064) );
  BUFx2_ASAP7_75t_R register___U7604 ( .A(register__n13333), .Y(register__n4065) );
  BUFx2_ASAP7_75t_R register___U7605 ( .A(register__n4067), .Y(register__n4066) );
  BUFx2_ASAP7_75t_R register___U7606 ( .A(register__n4071), .Y(register__n4070) );
  BUFx2_ASAP7_75t_R register___U7607 ( .A(register__n13090), .Y(register__n4071) );
  BUFx2_ASAP7_75t_R register___U7608 ( .A(register__n4073), .Y(register__n4072) );
  BUFx2_ASAP7_75t_R register___U7609 ( .A(register__n13108), .Y(register__n4073) );
  BUFx2_ASAP7_75t_R register___U7610 ( .A(register__n4075), .Y(register__n4074) );
  BUFx2_ASAP7_75t_R register___U7611 ( .A(register__n13100), .Y(register__n4075) );
  BUFx2_ASAP7_75t_R register___U7612 ( .A(register__n4077), .Y(register__n4076) );
  BUFx2_ASAP7_75t_R register___U7613 ( .A(register__n4079), .Y(register__n4078) );
  BUFx2_ASAP7_75t_R register___U7614 ( .A(register__n12880), .Y(register__n4079) );
  BUFx2_ASAP7_75t_R register___U7615 ( .A(register__n4081), .Y(register__n4080) );
  BUFx2_ASAP7_75t_R register___U7616 ( .A(register__n13201), .Y(register__n4081) );
  BUFx2_ASAP7_75t_R register___U7617 ( .A(register__n4089), .Y(register__n4088) );
  BUFx2_ASAP7_75t_R register___U7618 ( .A(register__n13106), .Y(register__n4089) );
  BUFx2_ASAP7_75t_R register___U7619 ( .A(register__n4091), .Y(register__n4090) );
  BUFx2_ASAP7_75t_R register___U7620 ( .A(register__n12984), .Y(register__n4091) );
  INVx6_ASAP7_75t_R register___U7621 ( .A(register__n12241), .Y(register__n12229) );
  BUFx2_ASAP7_75t_R register___U7622 ( .A(register__net135335), .Y(register__net135334) );
  BUFx2_ASAP7_75t_R register___U7623 ( .A(register__net35929), .Y(register__net135335) );
  BUFx2_ASAP7_75t_R register___U7624 ( .A(register__n4093), .Y(register__n4092) );
  BUFx2_ASAP7_75t_R register___U7625 ( .A(register__n13088), .Y(register__n4093) );
  BUFx2_ASAP7_75t_R register___U7626 ( .A(register__n4095), .Y(register__n4094) );
  BUFx2_ASAP7_75t_R register___U7627 ( .A(register__n13113), .Y(register__n4095) );
  BUFx3_ASAP7_75t_R register___U7628 ( .A(register__n4100), .Y(register__n4099) );
  BUFx2_ASAP7_75t_R register___U7629 ( .A(register__n11572), .Y(register__n4100) );
  BUFx3_ASAP7_75t_R register___U7630 ( .A(register__n4102), .Y(register__n4101) );
  BUFx2_ASAP7_75t_R register___U7631 ( .A(register__n11286), .Y(register__n4102) );
  BUFx2_ASAP7_75t_R register___U7632 ( .A(register__n6751), .Y(register__n4107) );
  BUFx3_ASAP7_75t_R register___U7633 ( .A(register__n4109), .Y(register__n4108) );
  BUFx2_ASAP7_75t_R register___U7634 ( .A(register__n10922), .Y(register__n4109) );
  BUFx2_ASAP7_75t_R register___U7635 ( .A(register__n5689), .Y(register__n4112) );
  BUFx3_ASAP7_75t_R register___U7636 ( .A(register__n4114), .Y(register__n4113) );
  BUFx2_ASAP7_75t_R register___U7637 ( .A(register__n10921), .Y(register__n4114) );
  BUFx3_ASAP7_75t_R register___U7638 ( .A(register__n4116), .Y(register__n4115) );
  BUFx2_ASAP7_75t_R register___U7639 ( .A(register__n11516), .Y(register__n4116) );
  BUFx12f_ASAP7_75t_R register___U7640 ( .A(register__net145201), .Y(register__net63210) );
  BUFx12f_ASAP7_75t_R register___U7641 ( .A(register__n2935), .Y(register__n11816) );
  BUFx12f_ASAP7_75t_R register___U7642 ( .A(register__net64984), .Y(register__net64980) );
  BUFx3_ASAP7_75t_R register___U7643 ( .A(register__net101209), .Y(register__net134932) );
  INVx1_ASAP7_75t_R register___U7644 ( .A(register__n2904), .Y(register__n4123) );
  BUFx3_ASAP7_75t_R register___U7645 ( .A(register__n4125), .Y(register__n4124) );
  BUFx2_ASAP7_75t_R register___U7646 ( .A(Reg_data[142]), .Y(register__n4125) );
  OA22x2_ASAP7_75t_R register___U7647 ( .A1(register__net63250), .A2(register__n1416), .B1(register__net90537), .B2(
        n1418), .Y(register__n12986) );
  OA22x2_ASAP7_75t_R register___U7648 ( .A1(register__net63340), .A2(register__n665), .B1(register__register__n6651), .B2(register__n81), 
        .Y(register__n12808) );
  INVx1_ASAP7_75t_R register___U7649 ( .A(register__n3587), .Y(register__n4126) );
  OA22x2_ASAP7_75t_R register___U7650 ( .A1(register__n12057), .A2(register__n1974), .B1(register__n9975), .B2(register__n11796), 
        .Y(register__n12910) );
  OA22x2_ASAP7_75t_R register___U7651 ( .A1(register__n12316), .A2(register__n956), .B1(register__n9644), .B2(register__n960), 
        .Y(register__n13020) );
  AND3x1_ASAP7_75t_R register___U7652 ( .A(register__n12515), .B(register__n6760), .C(register__n6761), .Y(register__n12521) );
  BUFx2_ASAP7_75t_R register___U7653 ( .A(register__n4131), .Y(register__n4130) );
  BUFx2_ASAP7_75t_R register___U7654 ( .A(register__n12776), .Y(register__n4131) );
  BUFx2_ASAP7_75t_R register___U7655 ( .A(register__n4133), .Y(register__n4132) );
  BUFx2_ASAP7_75t_R register___U7656 ( .A(register__n12992), .Y(register__n4133) );
  BUFx2_ASAP7_75t_R register___U7657 ( .A(register__n4135), .Y(register__n4134) );
  BUFx2_ASAP7_75t_R register___U7658 ( .A(register__n13006), .Y(register__n4135) );
  BUFx2_ASAP7_75t_R register___U7659 ( .A(register__n4137), .Y(register__n4136) );
  BUFx2_ASAP7_75t_R register___U7660 ( .A(register__n13216), .Y(register__n4137) );
  BUFx2_ASAP7_75t_R register___U7661 ( .A(register__n4139), .Y(register__n4138) );
  BUFx2_ASAP7_75t_R register___U7662 ( .A(register__n13235), .Y(register__n4139) );
  BUFx2_ASAP7_75t_R register___U7663 ( .A(register__n4147), .Y(register__n4146) );
  BUFx2_ASAP7_75t_R register___U7664 ( .A(register__n12982), .Y(register__n4147) );
  BUFx2_ASAP7_75t_R register___U7665 ( .A(register__n12754), .Y(register__n4151) );
  INVx6_ASAP7_75t_R register___U7666 ( .A(register__n12246), .Y(register__n12234) );
  BUFx3_ASAP7_75t_R register___U7667 ( .A(register__n4159), .Y(register__n4158) );
  BUFx2_ASAP7_75t_R register___U7668 ( .A(register__n10876), .Y(register__n4159) );
  BUFx3_ASAP7_75t_R register___U7669 ( .A(register__n10878), .Y(register__n4160) );
  BUFx2_ASAP7_75t_R register___U7670 ( .A(register__n5692), .Y(register__n4161) );
  BUFx3_ASAP7_75t_R register___U7671 ( .A(register__n4163), .Y(register__n4162) );
  BUFx2_ASAP7_75t_R register___U7672 ( .A(register__n10875), .Y(register__n4163) );
  BUFx3_ASAP7_75t_R register___U7673 ( .A(register__n4168), .Y(register__n4167) );
  BUFx2_ASAP7_75t_R register___U7674 ( .A(register__n11715), .Y(register__n4168) );
  BUFx3_ASAP7_75t_R register___U7675 ( .A(register__n4170), .Y(register__n4169) );
  BUFx2_ASAP7_75t_R register___U7676 ( .A(register__n11718), .Y(register__n4170) );
  BUFx2_ASAP7_75t_R register___U7677 ( .A(register__n7057), .Y(register__n4171) );
  BUFx3_ASAP7_75t_R register___U7678 ( .A(register__n4174), .Y(register__n4173) );
  BUFx2_ASAP7_75t_R register___U7679 ( .A(register__n11239), .Y(register__n4174) );
  BUFx3_ASAP7_75t_R register___U7680 ( .A(register__n4176), .Y(register__n4175) );
  BUFx2_ASAP7_75t_R register___U7681 ( .A(register__n11237), .Y(register__n4176) );
  AND4x1_ASAP7_75t_R register___U7682 ( .A(register__n455), .B(register__n11156), .C(register__n8250), .D(register__n11155), .Y(
        n8641) );
  AND4x1_ASAP7_75t_R register___U7683 ( .A(register__n8697), .B(register__n10907), .C(register__n10906), .D(register__n10908), 
        .Y(register__n7275) );
  AND4x1_ASAP7_75t_R register___U7684 ( .A(register__n10697), .B(register__n10698), .C(register__n10699), .D(register__n377), .Y(
        n7022) );
  BUFx3_ASAP7_75t_R register___U7685 ( .A(register__n8801), .Y(register__n4180) );
  BUFx4f_ASAP7_75t_R register___U7686 ( .A(register__n8801), .Y(register__n4181) );
  BUFx2_ASAP7_75t_R register___U7687 ( .A(register__n8801), .Y(register__n4182) );
  BUFx3_ASAP7_75t_R register___U7688 ( .A(register__net101199), .Y(register__net134033) );
  BUFx12f_ASAP7_75t_R register___U7689 ( .A(register__net89566), .Y(register__net89565) );
  OA22x2_ASAP7_75t_R register___U7690 ( .A1(register__net64664), .A2(register__n1416), .B1(register__n9786), .B2(register__n1418), 
        .Y(register__n13002) );
  OA22x2_ASAP7_75t_R register___U7691 ( .A1(register__n12289), .A2(register__n665), .B1(register__n8504), .B2(register__n81), .Y(
        n12812) );
  INVx1_ASAP7_75t_R register___U7692 ( .A(register__n2917), .Y(register__n4185) );
  OA22x2_ASAP7_75t_R register___U7693 ( .A1(register__net62988), .A2(register__n3337), .B1(register__n8169), .B2(register__n2856), 
        .Y(register__n13265) );
  INVx1_ASAP7_75t_R register___U7694 ( .A(register__n13265), .Y(register__n4186) );
  OA22x2_ASAP7_75t_R register___U7695 ( .A1(register__n12259), .A2(register__n337), .B1(register__n9625), .B2(register__n343), 
        .Y(register__n12729) );
  INVx1_ASAP7_75t_R register___U7696 ( .A(register__n3285), .Y(register__n4187) );
  OA22x2_ASAP7_75t_R register___U7697 ( .A1(register__net147310), .A2(register__n1973), .B1(register__net89997), .B2(
        n2892), .Y(register__n12912) );
  INVx1_ASAP7_75t_R register___U7698 ( .A(register__n2939), .Y(register__n4188) );
  OA22x2_ASAP7_75t_R register___U7699 ( .A1(register__net63166), .A2(register__n1415), .B1(register__net96903), .B2(
        n1418), .Y(register__n12985) );
  INVx1_ASAP7_75t_R register___U7700 ( .A(register__n3486), .Y(register__n4189) );
  OA22x2_ASAP7_75t_R register___U7701 ( .A1(register__n12056), .A2(register__n952), .B1(register__n9648), .B2(register__n960), 
        .Y(register__n13030) );
  OA22x2_ASAP7_75t_R register___U7702 ( .A1(register__net64840), .A2(register__n1755), .B1(register__net90789), .B2(
        n3821), .Y(register__n13142) );
  OA22x2_ASAP7_75t_R register___U7703 ( .A1(register__net63178), .A2(register__n11730), .B1(register__net88913), .B2(
        n1164), .Y(register__n13364) );
  INVx1_ASAP7_75t_R register___U7704 ( .A(register__n3160), .Y(register__n4190) );
  BUFx2_ASAP7_75t_R register___U7705 ( .A(register__n5986), .Y(register__n4191) );
  BUFx2_ASAP7_75t_R register___U7706 ( .A(register__n6398), .Y(register__n4192) );
  BUFx3_ASAP7_75t_R register___U7707 ( .A(register__n4196), .Y(register__n4195) );
  INVx6_ASAP7_75t_R register___U7708 ( .A(register__n12273), .Y(register__n12262) );
  BUFx12f_ASAP7_75t_R register___U7709 ( .A(register__n5034), .Y(register__n4197) );
  BUFx6f_ASAP7_75t_R register___U7710 ( .A(register__net64382), .Y(register__net133741) );
  BUFx12f_ASAP7_75t_R register___U7711 ( .A(register__net64382), .Y(register__net133742) );
  BUFx2_ASAP7_75t_R register___U7712 ( .A(register__n12799), .Y(register__n4205) );
  BUFx2_ASAP7_75t_R register___U7713 ( .A(register__n4211), .Y(register__n4210) );
  BUFx2_ASAP7_75t_R register___U7714 ( .A(register__n13249), .Y(register__n4211) );
  BUFx2_ASAP7_75t_R register___U7715 ( .A(register__n4215), .Y(register__n4214) );
  BUFx2_ASAP7_75t_R register___U7716 ( .A(register__n13082), .Y(register__n4215) );
  BUFx2_ASAP7_75t_R register___U7717 ( .A(register__n4217), .Y(register__n4216) );
  BUFx12f_ASAP7_75t_R register___U7718 ( .A(register__n12294), .Y(register__n12304) );
  BUFx3_ASAP7_75t_R register___U7719 ( .A(register__n4222), .Y(register__n4221) );
  BUFx2_ASAP7_75t_R register___U7720 ( .A(register__n11441), .Y(register__n4222) );
  BUFx2_ASAP7_75t_R register___U7721 ( .A(register__n6746), .Y(register__n4225) );
  BUFx3_ASAP7_75t_R register___U7722 ( .A(register__n4229), .Y(register__n4228) );
  BUFx2_ASAP7_75t_R register___U7723 ( .A(register__n11259), .Y(register__n4229) );
  BUFx3_ASAP7_75t_R register___U7724 ( .A(register__n4232), .Y(register__n4231) );
  BUFx2_ASAP7_75t_R register___U7725 ( .A(register__n11256), .Y(register__n4232) );
  BUFx3_ASAP7_75t_R register___U7726 ( .A(register__n4234), .Y(register__n4233) );
  BUFx2_ASAP7_75t_R register___U7727 ( .A(register__n11257), .Y(register__n4234) );
  BUFx3_ASAP7_75t_R register___U7728 ( .A(register__n4236), .Y(register__n4235) );
  BUFx2_ASAP7_75t_R register___U7729 ( .A(register__n11212), .Y(register__n4236) );
  BUFx3_ASAP7_75t_R register___U7730 ( .A(register__n4238), .Y(register__n4237) );
  BUFx2_ASAP7_75t_R register___U7731 ( .A(register__n11214), .Y(register__n4238) );
  BUFx2_ASAP7_75t_R register___U7732 ( .A(register__n7009), .Y(register__n4239) );
  BUFx3_ASAP7_75t_R register___U7733 ( .A(register__n4241), .Y(register__n4240) );
  BUFx2_ASAP7_75t_R register___U7734 ( .A(register__n11211), .Y(register__n4241) );
  BUFx2_ASAP7_75t_R register___U7735 ( .A(register__n5520), .Y(register__n4244) );
  BUFx2_ASAP7_75t_R register___U7736 ( .A(register__n7645), .Y(register__n4249) );
  BUFx3_ASAP7_75t_R register___U7737 ( .A(register__n4251), .Y(register__n4250) );
  BUFx2_ASAP7_75t_R register___U7738 ( .A(register__n10898), .Y(register__n4251) );
  BUFx3_ASAP7_75t_R register___U7739 ( .A(register__n4253), .Y(register__n4252) );
  BUFx2_ASAP7_75t_R register___U7740 ( .A(register__n11711), .Y(register__n4253) );
  BUFx3_ASAP7_75t_R register___U7741 ( .A(register__n4255), .Y(register__n4254) );
  BUFx2_ASAP7_75t_R register___U7742 ( .A(register__n11713), .Y(register__n4255) );
  BUFx3_ASAP7_75t_R register___U7743 ( .A(register__n4258), .Y(register__n4257) );
  BUFx2_ASAP7_75t_R register___U7744 ( .A(register__n11631), .Y(register__n4258) );
  BUFx3_ASAP7_75t_R register___U7745 ( .A(register__n4260), .Y(register__n4259) );
  BUFx2_ASAP7_75t_R register___U7746 ( .A(register__n11630), .Y(register__n4260) );
  BUFx12f_ASAP7_75t_R register___U7747 ( .A(register__n3044), .Y(register__n4266) );
  INVx6_ASAP7_75t_R register___U7748 ( .A(register__n4266), .Y(register__n12144) );
  BUFx3_ASAP7_75t_R register___U7749 ( .A(register__n4274), .Y(register__n4273) );
  BUFx2_ASAP7_75t_R register___U7750 ( .A(Reg_data[947]), .Y(register__n4274) );
  OA22x2_ASAP7_75t_R register___U7751 ( .A1(register__n12258), .A2(register__n2799), .B1(register__n6564), .B2(register__n3746), 
        .Y(register__n12813) );
  OA22x2_ASAP7_75t_R register___U7752 ( .A1(register__n12338), .A2(register__n2851), .B1(register__n10452), .B2(register__n3437), 
        .Y(register__n13270) );
  OA22x2_ASAP7_75t_R register___U7753 ( .A1(register__n12202), .A2(register__n337), .B1(register__n10487), .B2(register__n68), 
        .Y(register__n12731) );
  INVx1_ASAP7_75t_R register___U7754 ( .A(register__n3310), .Y(register__n4277) );
  OA22x2_ASAP7_75t_R register___U7755 ( .A1(register__net64848), .A2(register__n1914), .B1(register__net89993), .B2(
        n11784), .Y(register__n12913) );
  OA22x2_ASAP7_75t_R register___U7756 ( .A1(register__net64760), .A2(register__n953), .B1(register__net90905), .B2(register__n958), .Y(register__n13032) );
  OA22x2_ASAP7_75t_R register___U7757 ( .A1(register__net64924), .A2(register__n1755), .B1(register__n9690), .B2(register__n3821), 
        .Y(register__n13143) );
  INVx1_ASAP7_75t_R register___U7758 ( .A(register__n2913), .Y(register__n4279) );
  OA22x2_ASAP7_75t_R register___U7759 ( .A1(register__n12365), .A2(register__n11730), .B1(register__n10365), .B2(register__n1164), 
        .Y(register__n13367) );
  INVx1_ASAP7_75t_R register___U7760 ( .A(register__n3172), .Y(register__n4280) );
  BUFx2_ASAP7_75t_R register___U7761 ( .A(register__n6260), .Y(register__n4281) );
  INVx6_ASAP7_75t_R register___U7762 ( .A(register__net63212), .Y(register__net63176) );
  INVx6_ASAP7_75t_R register___U7763 ( .A(register__n3566), .Y(register__n11889) );
  INVx6_ASAP7_75t_R register___U7764 ( .A(register__net130019), .Y(register__net63244) );
  INVx4_ASAP7_75t_R register___U7765 ( .A(register__net145037), .Y(register__net109773) );
  BUFx3_ASAP7_75t_R register___U7766 ( .A(register__n4285), .Y(register__n4284) );
  BUFx2_ASAP7_75t_R register___U7767 ( .A(register__n11668), .Y(register__n4285) );
  BUFx3_ASAP7_75t_R register___U7768 ( .A(register__n4289), .Y(register__n4288) );
  BUFx2_ASAP7_75t_R register___U7769 ( .A(register__n11376), .Y(register__n4289) );
  BUFx12f_ASAP7_75t_R register___U7770 ( .A(register__net147289), .Y(register__net64470) );
  BUFx2_ASAP7_75t_R register___U7771 ( .A(register__n4294), .Y(register__n4293) );
  BUFx2_ASAP7_75t_R register___U7772 ( .A(register__n12674), .Y(register__n4294) );
  BUFx2_ASAP7_75t_R register___U7773 ( .A(register__n4301), .Y(register__n4300) );
  BUFx2_ASAP7_75t_R register___U7774 ( .A(register__n12681), .Y(register__n4301) );
  BUFx2_ASAP7_75t_R register___U7775 ( .A(register__n4303), .Y(register__n4302) );
  BUFx2_ASAP7_75t_R register___U7776 ( .A(register__n12539), .Y(register__n4303) );
  INVx1_ASAP7_75t_R register___U7777 ( .A(register__net62864), .Y(register__net132881) );
  BUFx12f_ASAP7_75t_R register___U7778 ( .A(register__net62848), .Y(register__net62864) );
  BUFx3_ASAP7_75t_R register___U7779 ( .A(register__n4307), .Y(register__n4306) );
  BUFx2_ASAP7_75t_R register___U7780 ( .A(register__n11549), .Y(register__n4307) );
  BUFx3_ASAP7_75t_R register___U7781 ( .A(register__n4311), .Y(register__n4310) );
  BUFx3_ASAP7_75t_R register___U7782 ( .A(register__n4313), .Y(register__n4312) );
  BUFx2_ASAP7_75t_R register___U7783 ( .A(register__n6414), .Y(register__n4314) );
  BUFx3_ASAP7_75t_R register___U7784 ( .A(register__n4316), .Y(register__n4315) );
  BUFx2_ASAP7_75t_R register___U7785 ( .A(register__n11532), .Y(register__n4316) );
  BUFx3_ASAP7_75t_R register___U7786 ( .A(register__n4318), .Y(register__n4317) );
  BUFx2_ASAP7_75t_R register___U7787 ( .A(register__n11292), .Y(register__n4318) );
  BUFx2_ASAP7_75t_R register___U7788 ( .A(register__n7264), .Y(register__n4319) );
  BUFx3_ASAP7_75t_R register___U7789 ( .A(register__n4321), .Y(register__n4320) );
  BUFx2_ASAP7_75t_R register___U7790 ( .A(register__n11289), .Y(register__n4321) );
  BUFx3_ASAP7_75t_R register___U7791 ( .A(register__n4323), .Y(register__n4322) );
  BUFx2_ASAP7_75t_R register___U7792 ( .A(register__n11233), .Y(register__n4323) );
  BUFx3_ASAP7_75t_R register___U7793 ( .A(register__n4325), .Y(register__n4324) );
  BUFx2_ASAP7_75t_R register___U7794 ( .A(register__n11232), .Y(register__n4325) );
  BUFx3_ASAP7_75t_R register___U7795 ( .A(register__n4327), .Y(register__n4326) );
  BUFx2_ASAP7_75t_R register___U7796 ( .A(register__n11235), .Y(register__n4327) );
  BUFx2_ASAP7_75t_R register___U7797 ( .A(register__n5699), .Y(register__n4328) );
  BUFx3_ASAP7_75t_R register___U7798 ( .A(register__n4330), .Y(register__n4329) );
  BUFx2_ASAP7_75t_R register___U7799 ( .A(register__n10626), .Y(register__n4330) );
  BUFx2_ASAP7_75t_R register___U7800 ( .A(register__n7643), .Y(register__n4333) );
  BUFx3_ASAP7_75t_R register___U7801 ( .A(register__n4341), .Y(register__n4340) );
  BUFx2_ASAP7_75t_R register___U7802 ( .A(register__n10648), .Y(register__n4341) );
  BUFx3_ASAP7_75t_R register___U7803 ( .A(register__n4343), .Y(register__n4342) );
  BUFx2_ASAP7_75t_R register___U7804 ( .A(register__n10989), .Y(register__n4343) );
  BUFx2_ASAP7_75t_R register___U7805 ( .A(register__n7311), .Y(register__n4344) );
  BUFx3_ASAP7_75t_R register___U7806 ( .A(register__n10986), .Y(register__n4347) );
  BUFx3_ASAP7_75t_R register___U7807 ( .A(register__n4349), .Y(register__n4348) );
  BUFx2_ASAP7_75t_R register___U7808 ( .A(register__n11461), .Y(register__n4349) );
  BUFx3_ASAP7_75t_R register___U7809 ( .A(register__n4351), .Y(register__n4350) );
  BUFx2_ASAP7_75t_R register___U7810 ( .A(register__n11463), .Y(register__n4351) );
  BUFx2_ASAP7_75t_R register___U7811 ( .A(register__n7015), .Y(register__n4352) );
  BUFx3_ASAP7_75t_R register___U7812 ( .A(register__n4354), .Y(register__n4353) );
  BUFx2_ASAP7_75t_R register___U7813 ( .A(register__n11673), .Y(register__n4354) );
  BUFx2_ASAP7_75t_R register___U7814 ( .A(register__n6421), .Y(register__n4355) );
  BUFx3_ASAP7_75t_R register___U7815 ( .A(register__n11671), .Y(register__n4356) );
  BUFx3_ASAP7_75t_R register___U7816 ( .A(register__n4360), .Y(register__n4359) );
  BUFx2_ASAP7_75t_R register___U7817 ( .A(register__n11627), .Y(register__n4360) );
  BUFx3_ASAP7_75t_R register___U7818 ( .A(register__n4362), .Y(register__n4361) );
  BUFx2_ASAP7_75t_R register___U7819 ( .A(register__n11218), .Y(register__n4362) );
  BUFx3_ASAP7_75t_R register___U7820 ( .A(register__n4364), .Y(register__n4363) );
  BUFx2_ASAP7_75t_R register___U7821 ( .A(register__n11215), .Y(register__n4364) );
  BUFx3_ASAP7_75t_R register___U7822 ( .A(register__n4366), .Y(register__n4365) );
  BUFx2_ASAP7_75t_R register___U7823 ( .A(register__n11216), .Y(register__n4366) );
  BUFx3_ASAP7_75t_R register___U7824 ( .A(register__n4368), .Y(register__n4367) );
  BUFx2_ASAP7_75t_R register___U7825 ( .A(register__n11402), .Y(register__n4368) );
  BUFx3_ASAP7_75t_R register___U7826 ( .A(register__n4370), .Y(register__n4369) );
  BUFx2_ASAP7_75t_R register___U7827 ( .A(register__n11405), .Y(register__n4370) );
  BUFx12f_ASAP7_75t_R register___U7828 ( .A(register__n2967), .Y(register__n4373) );
  BUFx3_ASAP7_75t_R register___U7829 ( .A(register__n4379), .Y(register__n4378) );
  BUFx2_ASAP7_75t_R register___U7830 ( .A(Reg_data[420]), .Y(register__n4379) );
  OA22x2_ASAP7_75t_R register___U7831 ( .A1(register__net63334), .A2(register__n101), .B1(register__n6654), .B2(register__n3302), 
        .Y(register__n12956) );
  INVx1_ASAP7_75t_R register___U7832 ( .A(register__n2973), .Y(register__n4381) );
  OA22x2_ASAP7_75t_R register___U7833 ( .A1(register__n12319), .A2(register__n1069), .B1(register__n82), .B2(register__n8799), 
        .Y(register__n12811) );
  OA22x2_ASAP7_75t_R register___U7834 ( .A1(register__net64770), .A2(register__n338), .B1(register__net90965), .B2(register__n342), .Y(register__n12741) );
  OA22x2_ASAP7_75t_R register___U7835 ( .A1(register__n12056), .A2(register__n1416), .B1(register__n10491), .B2(register__n1419), 
        .Y(register__n13001) );
  INVx1_ASAP7_75t_R register___U7836 ( .A(register__n3289), .Y(register__n4386) );
  OA22x2_ASAP7_75t_R register___U7837 ( .A1(register__net64844), .A2(register__n957), .B1(register__net90901), .B2(register__n960), .Y(register__n13033) );
  OA22x2_ASAP7_75t_R register___U7838 ( .A1(register__n11953), .A2(register__n1266), .B1(register__n10497), .B2(register__n3334), 
        .Y(register__n13146) );
  INVx1_ASAP7_75t_R register___U7839 ( .A(register__n13146), .Y(register__n4387) );
  OA22x2_ASAP7_75t_R register___U7840 ( .A1(register__n12310), .A2(register__n11730), .B1(register__n10367), .B2(register__n1164), 
        .Y(register__n13369) );
  INVx4_ASAP7_75t_R register___U7841 ( .A(register__n12012), .Y(register__n11997) );
  INVx6_ASAP7_75t_R register___U7842 ( .A(register__n12104), .Y(register__n12093) );
  BUFx2_ASAP7_75t_R register___U7843 ( .A(register__n4392), .Y(register__n4391) );
  BUFx2_ASAP7_75t_R register___U7844 ( .A(register__n12575), .Y(register__n4392) );
  INVx5_ASAP7_75t_R register___U7845 ( .A(register__net64890), .Y(register__net64860) );
  BUFx2_ASAP7_75t_R register___U7846 ( .A(register__n4400), .Y(register__n4399) );
  BUFx2_ASAP7_75t_R register___U7847 ( .A(register__n12631), .Y(register__n4400) );
  BUFx2_ASAP7_75t_R register___U7848 ( .A(register__n4402), .Y(register__n4401) );
  BUFx2_ASAP7_75t_R register___U7849 ( .A(register__n4404), .Y(register__n4403) );
  BUFx2_ASAP7_75t_R register___U7850 ( .A(register__n12646), .Y(register__n4404) );
  BUFx2_ASAP7_75t_R register___U7851 ( .A(register__n4408), .Y(register__n4407) );
  BUFx2_ASAP7_75t_R register___U7852 ( .A(register__n12665), .Y(register__n4408) );
  BUFx2_ASAP7_75t_R register___U7853 ( .A(register__n4410), .Y(register__n4409) );
  BUFx2_ASAP7_75t_R register___U7854 ( .A(register__n4416), .Y(register__n4415) );
  INVx6_ASAP7_75t_R register___U7855 ( .A(register__n4605), .Y(register__n12175) );
  BUFx2_ASAP7_75t_R register___U7856 ( .A(register__n4420), .Y(register__n4419) );
  BUFx2_ASAP7_75t_R register___U7857 ( .A(register__n13243), .Y(register__n4424) );
  BUFx2_ASAP7_75t_R register___U7858 ( .A(register__n7623), .Y(register__n4429) );
  BUFx2_ASAP7_75t_R register___U7859 ( .A(register__n12538), .Y(register__n4430) );
  BUFx3_ASAP7_75t_R register___U7860 ( .A(register__n4433), .Y(register__n4432) );
  BUFx2_ASAP7_75t_R register___U7861 ( .A(register__n11253), .Y(register__n4433) );
  BUFx3_ASAP7_75t_R register___U7862 ( .A(register__n4435), .Y(register__n4434) );
  BUFx2_ASAP7_75t_R register___U7863 ( .A(register__n11255), .Y(register__n4435) );
  BUFx2_ASAP7_75t_R register___U7864 ( .A(register__n5922), .Y(register__n4436) );
  BUFx3_ASAP7_75t_R register___U7865 ( .A(register__n4438), .Y(register__n4437) );
  BUFx2_ASAP7_75t_R register___U7866 ( .A(register__n11252), .Y(register__n4438) );
  BUFx3_ASAP7_75t_R register___U7867 ( .A(register__n4440), .Y(register__n4439) );
  BUFx2_ASAP7_75t_R register___U7868 ( .A(register__n11229), .Y(register__n4440) );
  BUFx3_ASAP7_75t_R register___U7869 ( .A(register__n10835), .Y(register__n4441) );
  BUFx2_ASAP7_75t_R register___U7870 ( .A(register__n6702), .Y(register__n4446) );
  BUFx3_ASAP7_75t_R register___U7871 ( .A(register__n4451), .Y(register__n4450) );
  BUFx2_ASAP7_75t_R register___U7872 ( .A(register__n10966), .Y(register__n4451) );
  BUFx2_ASAP7_75t_R register___U7873 ( .A(register__n10968), .Y(register__n4452) );
  BUFx2_ASAP7_75t_R register___U7874 ( .A(register__n6410), .Y(register__n4453) );
  BUFx3_ASAP7_75t_R register___U7875 ( .A(register__n4455), .Y(register__n4454) );
  BUFx2_ASAP7_75t_R register___U7876 ( .A(register__n10965), .Y(register__n4455) );
  BUFx3_ASAP7_75t_R register___U7877 ( .A(register__n10750), .Y(register__n4456) );
  BUFx2_ASAP7_75t_R register___U7878 ( .A(register__n6153), .Y(register__n4457) );
  BUFx3_ASAP7_75t_R register___U7879 ( .A(register__n4459), .Y(register__n4458) );
  BUFx2_ASAP7_75t_R register___U7880 ( .A(register__n10747), .Y(register__n4459) );
  BUFx3_ASAP7_75t_R register___U7881 ( .A(register__n4461), .Y(register__n4460) );
  BUFx2_ASAP7_75t_R register___U7882 ( .A(register__n11319), .Y(register__n4461) );
  BUFx3_ASAP7_75t_R register___U7883 ( .A(register__n4465), .Y(register__n4464) );
  BUFx2_ASAP7_75t_R register___U7884 ( .A(register__n11317), .Y(register__n4465) );
  BUFx3_ASAP7_75t_R register___U7885 ( .A(register__n4467), .Y(register__n4466) );
  BUFx2_ASAP7_75t_R register___U7886 ( .A(register__n11599), .Y(register__n4467) );
  BUFx3_ASAP7_75t_R register___U7887 ( .A(register__n4469), .Y(register__n4468) );
  BUFx2_ASAP7_75t_R register___U7888 ( .A(register__n11596), .Y(register__n4469) );
  BUFx3_ASAP7_75t_R register___U7889 ( .A(register__n4471), .Y(register__n4470) );
  OR2x2_ASAP7_75t_R register___U7890 ( .A(register__n4473), .B(register__n5899), .Y(register__n4472) );
  BUFx2_ASAP7_75t_R register___U7891 ( .A(register__n5898), .Y(register__n4473) );
  NOR2x1p5_ASAP7_75t_R register___U7892 ( .A(register__n10460), .B(register__n970), .Y(register__n5898) );
  NOR2x1p5_ASAP7_75t_R register___U7893 ( .A(register__n11952), .B(register__n985), .Y(register__n5899) );
  BUFx12f_ASAP7_75t_R register___U7894 ( .A(register__n11890), .Y(register__n4474) );
  BUFx12f_ASAP7_75t_R register___U7895 ( .A(register__n11740), .Y(register__n4475) );
  BUFx12f_ASAP7_75t_R register___U7896 ( .A(register__net131433), .Y(register__net64972) );
  BUFx3_ASAP7_75t_R register___U7897 ( .A(register__n4480), .Y(register__n4479) );
  BUFx2_ASAP7_75t_R register___U7898 ( .A(Reg_data[179]), .Y(register__n4480) );
  OA22x2_ASAP7_75t_R register___U7899 ( .A1(register__n11958), .A2(register__n2811), .B1(register__n6272), .B2(register__n2808), 
        .Y(register__n12886) );
  INVx1_ASAP7_75t_R register___U7900 ( .A(register__n12886), .Y(register__n4481) );
  INVx1_ASAP7_75t_R register___U7901 ( .A(register__n2946), .Y(register__n4483) );
  OA22x2_ASAP7_75t_R register___U7902 ( .A1(register__n12400), .A2(register__n100), .B1(register__n6964), .B2(register__n3185), 
        .Y(register__n12953) );
  INVx1_ASAP7_75t_R register___U7903 ( .A(register__n3080), .Y(register__n4484) );
  OA22x2_ASAP7_75t_R register___U7904 ( .A1(register__n12312), .A2(register__n1049), .B1(register__n10020), .B2(register__n3295), 
        .Y(register__n13271) );
  INVx1_ASAP7_75t_R register___U7905 ( .A(register__n13271), .Y(register__n4485) );
  OA22x2_ASAP7_75t_R register___U7906 ( .A1(register__net63172), .A2(register__n665), .B1(register__net90093), .B2(
        n3746), .Y(register__n12806) );
  INVx6_ASAP7_75t_R register___U7907 ( .A(register__net63206), .Y(register__net63172) );
  OA22x2_ASAP7_75t_R register___U7908 ( .A1(register__n12026), .A2(register__n1973), .B1(register__n9979), .B2(register__n11795), 
        .Y(register__n12915) );
  OA22x2_ASAP7_75t_R register___U7909 ( .A1(register__net64762), .A2(register__n1416), .B1(register__net90937), .B2(
        n1417), .Y(register__n13003) );
  INVx1_ASAP7_75t_R register___U7910 ( .A(register__n13003), .Y(register__n4487) );
  OA22x2_ASAP7_75t_R register___U7911 ( .A1(register__net64928), .A2(register__n953), .B1(register__n9650), .B2(register__n958), 
        .Y(register__n13034) );
  INVx1_ASAP7_75t_R register___U7912 ( .A(register__n3579), .Y(register__n4488) );
  OA22x2_ASAP7_75t_R register___U7913 ( .A1(register__n12254), .A2(register__n11730), .B1(register__n10369), .B2(register__n1164), 
        .Y(register__n13371) );
  INVx1_ASAP7_75t_R register___U7914 ( .A(register__n3222), .Y(register__n4489) );
  BUFx3_ASAP7_75t_R register___U7915 ( .A(register__n4492), .Y(register__n4491) );
  BUFx2_ASAP7_75t_R register___U7916 ( .A(register__n11534), .Y(register__n4492) );
  BUFx3_ASAP7_75t_R register___U7917 ( .A(register__n4494), .Y(register__n4493) );
  BUFx2_ASAP7_75t_R register___U7918 ( .A(register__n11422), .Y(register__n4494) );
  BUFx12f_ASAP7_75t_R register___U7919 ( .A(register__net97365), .Y(register__net131056) );
  BUFx12f_ASAP7_75t_R register___U7920 ( .A(register__net97365), .Y(register__net131057) );
  BUFx12f_ASAP7_75t_R register___U7921 ( .A(register__net97365), .Y(register__net131058) );
  BUFx12f_ASAP7_75t_R register___U7922 ( .A(register__net131058), .Y(register__net63200) );
  BUFx12f_ASAP7_75t_R register___U7923 ( .A(register__net132155), .Y(register__net63212) );
  BUFx12f_ASAP7_75t_R register___U7924 ( .A(register__net131057), .Y(register__net63208) );
  BUFx12f_ASAP7_75t_R register___U7925 ( .A(register__net131056), .Y(register__net63206) );
  BUFx12f_ASAP7_75t_R register___U7926 ( .A(register__net132155), .Y(register__net63202) );
  BUFx2_ASAP7_75t_R register___U7927 ( .A(register__n4496), .Y(register__n4495) );
  BUFx2_ASAP7_75t_R register___U7928 ( .A(register__n12727), .Y(register__n4496) );
  BUFx2_ASAP7_75t_R register___U7929 ( .A(register__n4500), .Y(register__n4499) );
  BUFx2_ASAP7_75t_R register___U7930 ( .A(register__n4502), .Y(register__n4501) );
  BUFx2_ASAP7_75t_R register___U7931 ( .A(register__n4504), .Y(register__n4503) );
  BUFx2_ASAP7_75t_R register___U7932 ( .A(register__n4508), .Y(register__n4507) );
  BUFx2_ASAP7_75t_R register___U7933 ( .A(register__n13327), .Y(register__n4508) );
  BUFx2_ASAP7_75t_R register___U7934 ( .A(register__n4510), .Y(register__n4509) );
  BUFx2_ASAP7_75t_R register___U7935 ( .A(register__n4512), .Y(register__n4511) );
  BUFx2_ASAP7_75t_R register___U7936 ( .A(register__n12615), .Y(register__n4512) );
  BUFx2_ASAP7_75t_R register___U7937 ( .A(register__n4514), .Y(register__n4513) );
  BUFx2_ASAP7_75t_R register___U7938 ( .A(register__n12632), .Y(register__n4514) );
  BUFx2_ASAP7_75t_R register___U7939 ( .A(register__n4516), .Y(register__n4515) );
  BUFx2_ASAP7_75t_R register___U7940 ( .A(register__n4520), .Y(register__n4519) );
  BUFx2_ASAP7_75t_R register___U7941 ( .A(register__n13236), .Y(register__n4520) );
  BUFx2_ASAP7_75t_R register___U7942 ( .A(register__n4526), .Y(register__n4525) );
  BUFx2_ASAP7_75t_R register___U7943 ( .A(register__n4530), .Y(register__n4529) );
  BUFx2_ASAP7_75t_R register___U7944 ( .A(register__n4532), .Y(register__n4531) );
  BUFx2_ASAP7_75t_R register___U7945 ( .A(register__n4534), .Y(register__n4533) );
  BUFx2_ASAP7_75t_R register___U7946 ( .A(register__n4536), .Y(register__n4535) );
  BUFx2_ASAP7_75t_R register___U7947 ( .A(register__n12722), .Y(register__n4536) );
  BUFx2_ASAP7_75t_R register___U7948 ( .A(register__n4538), .Y(register__n4537) );
  BUFx2_ASAP7_75t_R register___U7949 ( .A(register__n13221), .Y(register__n4538) );
  BUFx2_ASAP7_75t_R register___U7950 ( .A(register__n4540), .Y(register__n4539) );
  BUFx2_ASAP7_75t_R register___U7951 ( .A(register__n12748), .Y(register__n4540) );
  BUFx2_ASAP7_75t_R register___U7952 ( .A(register__n4544), .Y(register__n4543) );
  BUFx2_ASAP7_75t_R register___U7953 ( .A(register__n13310), .Y(register__n4544) );
  BUFx2_ASAP7_75t_R register___U7954 ( .A(register__n5375), .Y(register__n4545) );
  BUFx12f_ASAP7_75t_R register___U7955 ( .A(register__net142401), .Y(register__net130835) );
  BUFx3_ASAP7_75t_R register___U7956 ( .A(register__n4548), .Y(register__n4547) );
  BUFx2_ASAP7_75t_R register___U7957 ( .A(register__n11569), .Y(register__n4548) );
  BUFx3_ASAP7_75t_R register___U7958 ( .A(register__n4550), .Y(register__n4549) );
  BUFx2_ASAP7_75t_R register___U7959 ( .A(register__n11568), .Y(register__n4550) );
  BUFx2_ASAP7_75t_R register___U7960 ( .A(register__n5913), .Y(register__n4553) );
  BUFx3_ASAP7_75t_R register___U7961 ( .A(register__n4555), .Y(register__n4554) );
  BUFx2_ASAP7_75t_R register___U7962 ( .A(register__n10851), .Y(register__n4555) );
  BUFx3_ASAP7_75t_R register___U7963 ( .A(register__n11359), .Y(register__n4559) );
  BUFx3_ASAP7_75t_R register___U7964 ( .A(register__n4561), .Y(register__n4560) );
  BUFx2_ASAP7_75t_R register___U7965 ( .A(register__n11612), .Y(register__n4561) );
  BUFx2_ASAP7_75t_R register___U7966 ( .A(register__n6158), .Y(register__n4562) );
  BUFx3_ASAP7_75t_R register___U7967 ( .A(register__n4564), .Y(register__n4563) );
  BUFx3_ASAP7_75t_R register___U7968 ( .A(register__n11073), .Y(register__n4565) );
  BUFx3_ASAP7_75t_R register___U7969 ( .A(register__n4567), .Y(register__n4566) );
  BUFx2_ASAP7_75t_R register___U7970 ( .A(register__n11071), .Y(register__n4567) );
  BUFx2_ASAP7_75t_R register___U7971 ( .A(register__n11070), .Y(register__n4568) );
  BUFx2_ASAP7_75t_R register___U7972 ( .A(register__n7650), .Y(register__n4569) );
  BUFx3_ASAP7_75t_R register___U7973 ( .A(register__n4571), .Y(register__n4570) );
  BUFx2_ASAP7_75t_R register___U7974 ( .A(register__n11653), .Y(register__n4571) );
  BUFx2_ASAP7_75t_R register___U7975 ( .A(register__n7919), .Y(register__n4572) );
  BUFx3_ASAP7_75t_R register___U7976 ( .A(register__n4574), .Y(register__n4573) );
  BUFx2_ASAP7_75t_R register___U7977 ( .A(register__n11650), .Y(register__n4574) );
  BUFx3_ASAP7_75t_R register___U7978 ( .A(register__n4581), .Y(register__n4580) );
  BUFx2_ASAP7_75t_R register___U7979 ( .A(register__n11551), .Y(register__n4581) );
  CKINVDCx10_ASAP7_75t_R register___U7980 ( .A(register__net64718), .Y(register__net64684) );
  INVx1_ASAP7_75t_R register___U7981 ( .A(register__n3785), .Y(register__n4584) );
  OA22x2_ASAP7_75t_R register___U7982 ( .A1(register__n12121), .A2(register__n115), .B1(register__n10233), .B2(register__n1639), 
        .Y(register__n12764) );
  INVx1_ASAP7_75t_R register___U7983 ( .A(register__n12764), .Y(register__n4585) );
  OA22x2_ASAP7_75t_R register___U7984 ( .A1(register__n12174), .A2(register__n1643), .B1(register__n8490), .B2(register__n1628), 
        .Y(register__n12763) );
  OA22x2_ASAP7_75t_R register___U7985 ( .A1(register__net63258), .A2(register__n339), .B1(register__net109926), .B2(
        n345), .Y(register__n12723) );
  OA22x2_ASAP7_75t_R register___U7986 ( .A1(register__net62654), .A2(register__n577), .B1(register__n9130), .B2(register__n579), 
        .Y(register__n13208) );
  INVx1_ASAP7_75t_R register___U7987 ( .A(register__n13208), .Y(register__n4586) );
  OA22x2_ASAP7_75t_R register___U7988 ( .A1(register__n12177), .A2(register__n107), .B1(register__n7680), .B2(register__n1517), 
        .Y(register__n12594) );
  OA22x2_ASAP7_75t_R register___U7989 ( .A1(register__n12167), .A2(register__n2851), .B1(register__n10201), .B2(register__n3339), 
        .Y(register__n13275) );
  INVx1_ASAP7_75t_R register___U7990 ( .A(register__n13275), .Y(register__n4588) );
  OA22x2_ASAP7_75t_R register___U7991 ( .A1(register__n11994), .A2(register__n337), .B1(register__n9632), .B2(register__n345), 
        .Y(register__n12744) );
  INVx1_ASAP7_75t_R register___U7992 ( .A(register__n3762), .Y(register__n4589) );
  OA22x2_ASAP7_75t_R register___U7993 ( .A1(register__n12344), .A2(register__n1069), .B1(register__n9945), .B2(register__n81), 
        .Y(register__n12810) );
  INVx1_ASAP7_75t_R register___U7994 ( .A(register__n3193), .Y(register__n4590) );
  OA22x2_ASAP7_75t_R register___U7995 ( .A1(register__n11991), .A2(register__n1974), .B1(register__n9981), .B2(register__n11783), 
        .Y(register__n12916) );
  OA22x2_ASAP7_75t_R register___U7996 ( .A1(register__net64920), .A2(register__n1416), .B1(register__n8761), .B2(register__n1417), 
        .Y(register__n13005) );
  INVx1_ASAP7_75t_R register___U7997 ( .A(register__n3398), .Y(register__n4591) );
  OA22x2_ASAP7_75t_R register___U7998 ( .A1(register__n3441), .A2(register__n957), .B1(register__n9652), .B2(register__n959), .Y(
        n13035) );
  OA22x2_ASAP7_75t_R register___U7999 ( .A1(register__n12051), .A2(register__n11730), .B1(register__n10371), .B2(register__n1164), 
        .Y(register__n13381) );
  INVx1_ASAP7_75t_R register___U8000 ( .A(register__n3269), .Y(register__n4592) );
  OA22x2_ASAP7_75t_R register___U8001 ( .A1(register__n12146), .A2(register__n1755), .B1(register__n9718), .B2(register__n3821), 
        .Y(register__n13134) );
  OA22x2_ASAP7_75t_R register___U8002 ( .A1(register__n12317), .A2(register__n100), .B1(register__n9278), .B2(register__n11770), 
        .Y(register__n12959) );
  INVx1_ASAP7_75t_R register___U8003 ( .A(register__n2879), .Y(register__n4594) );
  BUFx12f_ASAP7_75t_R register___U8004 ( .A(register__n12049), .Y(register__n4595) );
  BUFx12f_ASAP7_75t_R register___U8005 ( .A(register__n3320), .Y(register__n12216) );
  BUFx12f_ASAP7_75t_R register___U8006 ( .A(register__C6422_net69812), .Y(register__net130087) );
  INVx1_ASAP7_75t_R register___U8007 ( .A(register__n12352), .Y(register__n4596) );
  BUFx6f_ASAP7_75t_R register___U8008 ( .A(register__n5346), .Y(register__n12352) );
  BUFx12f_ASAP7_75t_R register___U8009 ( .A(register__net139893), .Y(register__net130019) );
  BUFx12f_ASAP7_75t_R register___U8010 ( .A(register__net139892), .Y(register__net130020) );
  BUFx2_ASAP7_75t_R register___U8011 ( .A(register__n4598), .Y(register__n4597) );
  BUFx2_ASAP7_75t_R register___U8012 ( .A(register__n12572), .Y(register__n4598) );
  BUFx2_ASAP7_75t_R register___U8013 ( .A(register__n4600), .Y(register__n4599) );
  BUFx2_ASAP7_75t_R register___U8014 ( .A(register__n12555), .Y(register__n4600) );
  BUFx12f_ASAP7_75t_R register___U8015 ( .A(register__n4606), .Y(register__n4605) );
  BUFx12f_ASAP7_75t_R register___U8016 ( .A(register__n3599), .Y(register__n4606) );
  BUFx12f_ASAP7_75t_R register___U8017 ( .A(register__n4747), .Y(register__n12188) );
  BUFx12f_ASAP7_75t_R register___U8018 ( .A(register__n3597), .Y(register__n12330) );
  BUFx12f_ASAP7_75t_R register___U8019 ( .A(register__net120674), .Y(register__net129901) );
  BUFx6f_ASAP7_75t_R register___U8020 ( .A(register__net129901), .Y(register__net64050) );
  BUFx12f_ASAP7_75t_R register___U8021 ( .A(register__net129901), .Y(register__net64044) );
  BUFx3_ASAP7_75t_R register___U8022 ( .A(register__n4611), .Y(register__n4610) );
  BUFx2_ASAP7_75t_R register___U8023 ( .A(register__n11248), .Y(register__n4611) );
  BUFx3_ASAP7_75t_R register___U8024 ( .A(register__n4613), .Y(register__n4612) );
  BUFx2_ASAP7_75t_R register___U8025 ( .A(register__n11163), .Y(register__n4613) );
  BUFx3_ASAP7_75t_R register___U8026 ( .A(register__n4615), .Y(register__n4614) );
  BUFx2_ASAP7_75t_R register___U8027 ( .A(register__n11162), .Y(register__n4615) );
  BUFx3_ASAP7_75t_R register___U8028 ( .A(register__n11010), .Y(register__n4618) );
  BUFx3_ASAP7_75t_R register___U8029 ( .A(register__n4620), .Y(register__n4619) );
  BUFx2_ASAP7_75t_R register___U8030 ( .A(register__n11009), .Y(register__n4620) );
  BUFx2_ASAP7_75t_R register___U8031 ( .A(register__n7909), .Y(register__n4621) );
  BUFx3_ASAP7_75t_R register___U8032 ( .A(register__n4626), .Y(register__n4625) );
  BUFx2_ASAP7_75t_R register___U8033 ( .A(register__n11689), .Y(register__n4626) );
  BUFx3_ASAP7_75t_R register___U8034 ( .A(register__n4628), .Y(register__n4627) );
  BUFx2_ASAP7_75t_R register___U8035 ( .A(register__n11589), .Y(register__n4628) );
  BUFx3_ASAP7_75t_R register___U8036 ( .A(register__n4630), .Y(register__n4629) );
  BUFx2_ASAP7_75t_R register___U8037 ( .A(register__n11588), .Y(register__n4630) );
  BUFx12f_ASAP7_75t_R register___U8038 ( .A(register__n3258), .Y(register__n4631) );
  BUFx12f_ASAP7_75t_R register___U8039 ( .A(register__net129693), .Y(register__net129691) );
  BUFx12f_ASAP7_75t_R register___U8040 ( .A(register__net143812), .Y(register__net63042) );
  BUFx12f_ASAP7_75t_R register___U8041 ( .A(register__net63052), .Y(register__net63048) );
  BUFx12f_ASAP7_75t_R register___U8042 ( .A(register__n4638), .Y(register__n4637) );
  BUFx12f_ASAP7_75t_R register___U8043 ( .A(register__n11867), .Y(register__n4638) );
  BUFx12f_ASAP7_75t_R register___U8044 ( .A(register__n3416), .Y(register__n11867) );
  BUFx12f_ASAP7_75t_R register___U8045 ( .A(register__net73059), .Y(register__net73055) );
  BUFx12f_ASAP7_75t_R register___U8046 ( .A(register__net134981), .Y(register__net64958) );
  BUFx12f_ASAP7_75t_R register___U8047 ( .A(register__n2986), .Y(register__n12161) );
  BUFx12f_ASAP7_75t_R register___U8048 ( .A(register__n4639), .Y(register__n12155) );
  BUFx12f_ASAP7_75t_R register___U8049 ( .A(register__n3513), .Y(register__n12163) );
  INVx1_ASAP7_75t_R register___U8050 ( .A(register__n3613), .Y(register__n4642) );
  OA22x2_ASAP7_75t_R register___U8051 ( .A1(register__net63180), .A2(register__n1961), .B1(register__net106940), .B2(
        n1525), .Y(register__n12584) );
  INVx1_ASAP7_75t_R register___U8052 ( .A(register__n3428), .Y(register__n4643) );
  OA22x2_ASAP7_75t_R register___U8053 ( .A1(register__n12059), .A2(register__n665), .B1(register__n8785), .B2(register__n81), .Y(
        n12823) );
  INVx1_ASAP7_75t_R register___U8054 ( .A(register__n3287), .Y(register__n4644) );
  OA22x2_ASAP7_75t_R register___U8055 ( .A1(register__n11957), .A2(register__n1973), .B1(register__n9983), .B2(register__n11789), 
        .Y(register__n12917) );
  OA22x2_ASAP7_75t_R register___U8056 ( .A1(register__n11989), .A2(register__n953), .B1(register__n9654), .B2(register__n960), 
        .Y(register__n13036) );
  OA22x2_ASAP7_75t_R register___U8057 ( .A1(register__net63156), .A2(register__n11868), .B1(register__net89889), .B2(
        n11748), .Y(register__n13267) );
  OA22x2_ASAP7_75t_R register___U8058 ( .A1(register__net64832), .A2(register__n11730), .B1(register__net88889), .B2(
        n1164), .Y(register__n13383) );
  INVx1_ASAP7_75t_R register___U8059 ( .A(register__n3291), .Y(register__n4646) );
  OA22x2_ASAP7_75t_R register___U8060 ( .A1(register__net64350), .A2(register__n336), .B1(register__net90681), .B2(register__n68), 
        .Y(register__n12736) );
  OA22x2_ASAP7_75t_R register___U8061 ( .A1(register__n3411), .A2(register__n100), .B1(register__n9280), .B2(register__n11768), 
        .Y(register__n12961) );
  OA22x2_ASAP7_75t_R register___U8062 ( .A1(register__n12406), .A2(register__n1755), .B1(register__n9766), .B2(register__n3334), 
        .Y(register__n13121) );
  BUFx12f_ASAP7_75t_R register___U8063 ( .A(register__n6404), .Y(register__n4650) );
  INVx5_ASAP7_75t_R register___U8064 ( .A(register__n11978), .Y(register__n11961) );
  INVx6_ASAP7_75t_R register___U8065 ( .A(register__n12333), .Y(register__n12321) );
  BUFx2_ASAP7_75t_R register___U8066 ( .A(register__n4652), .Y(register__n4651) );
  BUFx2_ASAP7_75t_R register___U8067 ( .A(register__n4654), .Y(register__n4653) );
  BUFx2_ASAP7_75t_R register___U8068 ( .A(register__n13067), .Y(register__n4654) );
  BUFx2_ASAP7_75t_R register___U8069 ( .A(register__n4656), .Y(register__n4655) );
  BUFx2_ASAP7_75t_R register___U8070 ( .A(register__n13294), .Y(register__n4656) );
  BUFx2_ASAP7_75t_R register___U8071 ( .A(register__n12707), .Y(register__n4658) );
  BUFx2_ASAP7_75t_R register___U8072 ( .A(register__n12705), .Y(register__n4660) );
  BUFx2_ASAP7_75t_R register___U8073 ( .A(register__n4664), .Y(register__n4663) );
  BUFx2_ASAP7_75t_R register___U8074 ( .A(register__n4666), .Y(register__n4665) );
  BUFx2_ASAP7_75t_R register___U8075 ( .A(register__n4668), .Y(register__n4667) );
  BUFx2_ASAP7_75t_R register___U8076 ( .A(register__n4670), .Y(register__n4669) );
  BUFx2_ASAP7_75t_R register___U8077 ( .A(register__n4672), .Y(register__n4671) );
  BUFx2_ASAP7_75t_R register___U8078 ( .A(register__n12683), .Y(register__n4672) );
  BUFx2_ASAP7_75t_R register___U8079 ( .A(register__n4676), .Y(register__n4675) );
  BUFx3_ASAP7_75t_R register___U8080 ( .A(register__n4685), .Y(register__n4684) );
  BUFx2_ASAP7_75t_R register___U8081 ( .A(register__n11207), .Y(register__n4685) );
  BUFx3_ASAP7_75t_R register___U8082 ( .A(register__n4687), .Y(register__n4686) );
  BUFx2_ASAP7_75t_R register___U8083 ( .A(register__n11208), .Y(register__n4687) );
  BUFx3_ASAP7_75t_R register___U8084 ( .A(register__n4689), .Y(register__n4688) );
  BUFx2_ASAP7_75t_R register___U8085 ( .A(register__n10926), .Y(register__n4689) );
  BUFx3_ASAP7_75t_R register___U8086 ( .A(register__n4691), .Y(register__n4690) );
  BUFx2_ASAP7_75t_R register___U8087 ( .A(register__n10925), .Y(register__n4691) );
  BUFx3_ASAP7_75t_R register___U8088 ( .A(register__n4693), .Y(register__n4692) );
  BUFx2_ASAP7_75t_R register___U8089 ( .A(register__n10927), .Y(register__n4693) );
  BUFx3_ASAP7_75t_R register___U8090 ( .A(register__n4695), .Y(register__n4694) );
  BUFx2_ASAP7_75t_R register___U8091 ( .A(register__n11398), .Y(register__n4695) );
  BUFx3_ASAP7_75t_R register___U8092 ( .A(register__n4697), .Y(register__n4696) );
  BUFx2_ASAP7_75t_R register___U8093 ( .A(register__n11399), .Y(register__n4697) );
  BUFx3_ASAP7_75t_R register___U8094 ( .A(register__n11357), .Y(register__n4701) );
  BUFx3_ASAP7_75t_R register___U8095 ( .A(register__n4709), .Y(register__n4708) );
  BUFx2_ASAP7_75t_R register___U8096 ( .A(register__n11026), .Y(register__n4709) );
  BUFx3_ASAP7_75t_R register___U8097 ( .A(register__n4711), .Y(register__n4710) );
  BUFx2_ASAP7_75t_R register___U8098 ( .A(register__n11029), .Y(register__n4711) );
  BUFx2_ASAP7_75t_R register___U8099 ( .A(register__n6427), .Y(register__n4712) );
  BUFx3_ASAP7_75t_R register___U8100 ( .A(register__n4714), .Y(register__n4713) );
  BUFx2_ASAP7_75t_R register___U8101 ( .A(register__n11089), .Y(register__n4714) );
  BUFx3_ASAP7_75t_R register___U8102 ( .A(register__n11090), .Y(register__n4715) );
  BUFx3_ASAP7_75t_R register___U8103 ( .A(register__n4719), .Y(register__n4718) );
  BUFx2_ASAP7_75t_R register___U8104 ( .A(register__n11595), .Y(register__n4719) );
  BUFx3_ASAP7_75t_R register___U8105 ( .A(register__n4722), .Y(register__n4721) );
  BUFx2_ASAP7_75t_R register___U8106 ( .A(register__n11375), .Y(register__n4722) );
  BUFx12f_ASAP7_75t_R register___U8107 ( .A(register__net141985), .Y(register__net62686) );
  AO22x1_ASAP7_75t_R register___U8108 ( .A1(register__n10493), .A2(register__n1867), .B1(register__n7994), .B2(register__n1354), 
        .Y(register__n10669) );
  BUFx3_ASAP7_75t_R register___U8109 ( .A(register__n4724), .Y(register__n4723) );
  BUFx2_ASAP7_75t_R register___U8110 ( .A(register__n10646), .Y(register__n4724) );
  BUFx3_ASAP7_75t_R register___U8111 ( .A(register__n4726), .Y(register__n4725) );
  BUFx2_ASAP7_75t_R register___U8112 ( .A(register__n10645), .Y(register__n4726) );
  BUFx12f_ASAP7_75t_R register___U8113 ( .A(register__n1326), .Y(register__n12413) );
  BUFx3_ASAP7_75t_R register___U8114 ( .A(register__n4731), .Y(register__n4730) );
  BUFx2_ASAP7_75t_R register___U8115 ( .A(register__n11606), .Y(register__n4731) );
  BUFx3_ASAP7_75t_R register___U8116 ( .A(register__n4733), .Y(register__n4732) );
  BUFx2_ASAP7_75t_R register___U8117 ( .A(register__n11607), .Y(register__n4733) );
  BUFx3_ASAP7_75t_R register___U8118 ( .A(register__n4735), .Y(register__n4734) );
  BUFx3_ASAP7_75t_R register___U8119 ( .A(register__n4737), .Y(register__n4736) );
  BUFx2_ASAP7_75t_R register___U8120 ( .A(register__n11712), .Y(register__n4737) );
  INVx1_ASAP7_75t_R register___U8121 ( .A(register__n11646), .Y(register__n4740) );
  BUFx3_ASAP7_75t_R register___U8122 ( .A(register__n4742), .Y(register__n4741) );
  BUFx2_ASAP7_75t_R register___U8123 ( .A(register__n11647), .Y(register__n4742) );
  BUFx3_ASAP7_75t_R register___U8124 ( .A(register__n4744), .Y(register__n4743) );
  BUFx2_ASAP7_75t_R register___U8125 ( .A(register__n11418), .Y(register__n4744) );
  BUFx12f_ASAP7_75t_R register___U8126 ( .A(register__n5043), .Y(register__n4747) );
  BUFx12f_ASAP7_75t_R register___U8127 ( .A(register__n12189), .Y(register__n4748) );
  BUFx3_ASAP7_75t_R register___U8128 ( .A(register__n4750), .Y(register__n4749) );
  BUFx2_ASAP7_75t_R register___U8129 ( .A(register__n10594), .Y(register__n4750) );
  BUFx3_ASAP7_75t_R register___U8130 ( .A(register__n4752), .Y(register__n4751) );
  BUFx2_ASAP7_75t_R register___U8131 ( .A(register__n10593), .Y(register__n4752) );
  BUFx2_ASAP7_75t_R register___U8132 ( .A(register__n8696), .Y(register__n4755) );
  BUFx3_ASAP7_75t_R register___U8133 ( .A(register__n9943), .Y(register__n4756) );
  BUFx4f_ASAP7_75t_R register___U8134 ( .A(register__n9943), .Y(register__n4757) );
  BUFx2_ASAP7_75t_R register___U8135 ( .A(register__n9943), .Y(register__n4758) );
  BUFx12f_ASAP7_75t_R register___U8136 ( .A(register__n1901), .Y(register__n11738) );
  INVx1_ASAP7_75t_R register___U8137 ( .A(register__n2841), .Y(register__n4759) );
  INVx1_ASAP7_75t_R register___U8138 ( .A(register__n3058), .Y(register__n4760) );
  INVx1_ASAP7_75t_R register___U8139 ( .A(register__n3061), .Y(register__n4761) );
  OA22x2_ASAP7_75t_R register___U8140 ( .A1(register__net63002), .A2(register__n2983), .B1(register__n7718), .B2(register__n12498), .Y(register__n12862) );
  INVx1_ASAP7_75t_R register___U8141 ( .A(register__n3661), .Y(register__n4762) );
  OA22x2_ASAP7_75t_R register___U8142 ( .A1(register__net62992), .A2(register__n1139), .B1(register__n7721), .B2(register__n1146), 
        .Y(register__n13152) );
  OA22x2_ASAP7_75t_R register___U8143 ( .A1(register__n12349), .A2(register__n113), .B1(register__n10479), .B2(register__n1524), 
        .Y(register__n12587) );
  INVx1_ASAP7_75t_R register___U8144 ( .A(register__n3458), .Y(register__n4763) );
  OA22x2_ASAP7_75t_R register___U8145 ( .A1(register__net63174), .A2(register__n1792), .B1(register__net90169), .B2(
        n1626), .Y(register__n12752) );
  INVx1_ASAP7_75t_R register___U8146 ( .A(register__n12752), .Y(register__n4764) );
  OA22x2_ASAP7_75t_R register___U8147 ( .A1(register__net64768), .A2(register__n665), .B1(register__net90081), .B2(register__n81), 
        .Y(register__n12825) );
  INVx1_ASAP7_75t_R register___U8148 ( .A(register__n3312), .Y(register__n4765) );
  OA22x2_ASAP7_75t_R register___U8149 ( .A1(register__n11928), .A2(register__n1973), .B1(register__n9985), .B2(register__n11797), 
        .Y(register__n12918) );
  INVx1_ASAP7_75t_R register___U8150 ( .A(register__n2954), .Y(register__n4766) );
  OA22x2_ASAP7_75t_R register___U8151 ( .A1(register__n11955), .A2(register__n955), .B1(register__n9656), .B2(register__n959), 
        .Y(register__n13037) );
  OA22x2_ASAP7_75t_R register___U8152 ( .A1(register__n12313), .A2(register__n578), .B1(register__n10056), .B2(register__n588), 
        .Y(register__n13218) );
  INVx1_ASAP7_75t_R register___U8153 ( .A(register__n4515), .Y(register__n4767) );
  OA22x2_ASAP7_75t_R register___U8154 ( .A1(register__net64328), .A2(register__n3719), .B1(register__net88885), .B2(
        n11848), .Y(register__n13378) );
  INVx1_ASAP7_75t_R register___U8155 ( .A(register__n13378), .Y(register__n4768) );
  OA22x2_ASAP7_75t_R register___U8156 ( .A1(register__n12149), .A2(register__n1412), .B1(register__n9746), .B2(register__n1417), 
        .Y(register__n12997) );
  OA22x2_ASAP7_75t_R register___U8157 ( .A1(register__n12149), .A2(register__n101), .B1(register__n9282), .B2(register__n11776), 
        .Y(register__n12966) );
  INVx6_ASAP7_75t_R register___U8158 ( .A(register__n12160), .Y(register__n12149) );
  BUFx2_ASAP7_75t_R register___U8159 ( .A(register__n8228), .Y(register__n4772) );
  BUFx2_ASAP7_75t_R register___U8160 ( .A(register__n4774), .Y(register__n4773) );
  BUFx2_ASAP7_75t_R register___U8161 ( .A(register__n12933), .Y(register__n4774) );
  BUFx2_ASAP7_75t_R register___U8162 ( .A(register__n4780), .Y(register__n4779) );
  BUFx2_ASAP7_75t_R register___U8163 ( .A(register__n12942), .Y(register__n4780) );
  BUFx6f_ASAP7_75t_R register___U8164 ( .A(register__n4727), .Y(register__n12414) );
  BUFx3_ASAP7_75t_R register___U8165 ( .A(register__n4788), .Y(register__n4787) );
  BUFx2_ASAP7_75t_R register___U8166 ( .A(register__n10970), .Y(register__n4788) );
  BUFx3_ASAP7_75t_R register___U8167 ( .A(register__n4790), .Y(register__n4789) );
  BUFx2_ASAP7_75t_R register___U8168 ( .A(register__n10969), .Y(register__n4790) );
  BUFx3_ASAP7_75t_R register___U8169 ( .A(register__n4792), .Y(register__n4791) );
  BUFx2_ASAP7_75t_R register___U8170 ( .A(register__n10971), .Y(register__n4792) );
  BUFx3_ASAP7_75t_R register___U8171 ( .A(register__n10774), .Y(register__n4793) );
  BUFx2_ASAP7_75t_R register___U8172 ( .A(register__n6716), .Y(register__n4794) );
  BUFx3_ASAP7_75t_R register___U8173 ( .A(register__n4796), .Y(register__n4795) );
  BUFx2_ASAP7_75t_R register___U8174 ( .A(register__n10772), .Y(register__n4796) );
  BUFx3_ASAP7_75t_R register___U8175 ( .A(register__n4798), .Y(register__n4797) );
  BUFx2_ASAP7_75t_R register___U8176 ( .A(register__n10712), .Y(register__n4798) );
  BUFx3_ASAP7_75t_R register___U8177 ( .A(register__n4800), .Y(register__n4799) );
  BUFx2_ASAP7_75t_R register___U8178 ( .A(register__n10815), .Y(register__n4800) );
  BUFx3_ASAP7_75t_R register___U8179 ( .A(register__n4802), .Y(register__n4801) );
  BUFx2_ASAP7_75t_R register___U8180 ( .A(register__n10992), .Y(register__n4802) );
  BUFx3_ASAP7_75t_R register___U8181 ( .A(register__n4804), .Y(register__n4803) );
  BUFx2_ASAP7_75t_R register___U8182 ( .A(register__n10990), .Y(register__n4804) );
  BUFx3_ASAP7_75t_R register___U8183 ( .A(register__n4806), .Y(register__n4805) );
  BUFx2_ASAP7_75t_R register___U8184 ( .A(register__n10991), .Y(register__n4806) );
  BUFx3_ASAP7_75t_R register___U8185 ( .A(register__n4808), .Y(register__n4807) );
  BUFx2_ASAP7_75t_R register___U8186 ( .A(register__n10794), .Y(register__n4808) );
  BUFx3_ASAP7_75t_R register___U8187 ( .A(register__n4810), .Y(register__n4809) );
  BUFx2_ASAP7_75t_R register___U8188 ( .A(register__n6707), .Y(register__n4811) );
  BUFx3_ASAP7_75t_R register___U8189 ( .A(register__n4814), .Y(register__n4813) );
  BUFx2_ASAP7_75t_R register___U8190 ( .A(register__n11048), .Y(register__n4814) );
  BUFx12f_ASAP7_75t_R register___U8191 ( .A(register__n3355), .Y(register__n4815) );
  BUFx12f_ASAP7_75t_R register___U8192 ( .A(register__n11914), .Y(register__n4818) );
  BUFx12f_ASAP7_75t_R register___U8193 ( .A(register__n3706), .Y(register__n11914) );
  BUFx12f_ASAP7_75t_R register___U8194 ( .A(register__net64788), .Y(register__net127693) );
  BUFx4f_ASAP7_75t_R register___U8195 ( .A(register__net136247), .Y(register__net64792) );
  BUFx6f_ASAP7_75t_R register___U8196 ( .A(register__net136248), .Y(register__net64794) );
  BUFx3_ASAP7_75t_R register___U8197 ( .A(register__n4821), .Y(register__n4820) );
  BUFx2_ASAP7_75t_R register___U8198 ( .A(register__n11138), .Y(register__n4821) );
  AND4x1_ASAP7_75t_R register___U8199 ( .A(register__n2053), .B(register__n4375), .C(register__n12519), .D(register__n12518), .Y(
        n12520) );
  BUFx3_ASAP7_75t_R register___U8200 ( .A(register__n4825), .Y(register__n4824) );
  BUFx2_ASAP7_75t_R register___U8201 ( .A(register__n10617), .Y(register__n4825) );
  BUFx3_ASAP7_75t_R register___U8202 ( .A(register__n4827), .Y(register__n4826) );
  BUFx2_ASAP7_75t_R register___U8203 ( .A(register__n10616), .Y(register__n4827) );
  BUFx2_ASAP7_75t_R register___U8204 ( .A(register__n8308), .Y(register__n4828) );
  BUFx3_ASAP7_75t_R register___U8205 ( .A(register__n4830), .Y(register__n4829) );
  BUFx2_ASAP7_75t_R register___U8206 ( .A(register__n10720), .Y(register__n4830) );
  BUFx3_ASAP7_75t_R register___U8207 ( .A(register__n4832), .Y(register__n4831) );
  BUFx2_ASAP7_75t_R register___U8208 ( .A(register__n10719), .Y(register__n4832) );
  BUFx12f_ASAP7_75t_R register___U8209 ( .A(register__n3701), .Y(register__n4834) );
  BUFx12f_ASAP7_75t_R register___U8210 ( .A(register__n3702), .Y(register__n4835) );
  BUFx12f_ASAP7_75t_R register___U8211 ( .A(register__n4835), .Y(register__n12333) );
  BUFx6f_ASAP7_75t_R register___U8212 ( .A(register__n4834), .Y(register__n12332) );
  BUFx12f_ASAP7_75t_R register___U8213 ( .A(register__n4839), .Y(register__n4838) );
  BUFx12f_ASAP7_75t_R register___U8214 ( .A(register__n5516), .Y(register__n11875) );
  BUFx12f_ASAP7_75t_R register___U8215 ( .A(register__net137521), .Y(register__net99879) );
  INVx6_ASAP7_75t_R register___U8216 ( .A(register__net99879), .Y(register__net127380) );
  BUFx12f_ASAP7_75t_R register___U8217 ( .A(register__n4845), .Y(register__n4844) );
  BUFx12f_ASAP7_75t_R register___U8218 ( .A(register__n3360), .Y(register__n4845) );
  CKINVDCx5p33_ASAP7_75t_R register___U8219 ( .A(register__net64684), .Y(register__net127351) );
  BUFx4f_ASAP7_75t_R register___U8220 ( .A(register__net127351), .Y(register__net64706) );
  BUFx3_ASAP7_75t_R register___U8221 ( .A(register__net127332), .Y(register__net127331) );
  BUFx2_ASAP7_75t_R register___U8222 ( .A(Reg_data[523]), .Y(register__net127332) );
  BUFx3_ASAP7_75t_R register___U8223 ( .A(register__net127328), .Y(register__net127327) );
  BUFx2_ASAP7_75t_R register___U8224 ( .A(Reg_data[906]), .Y(register__net127328) );
  OA22x2_ASAP7_75t_R register___U8225 ( .A1(register__net62648), .A2(register__n11730), .B1(register__n10415), .B2(
        n1164), .Y(register__n13358) );
  INVx1_ASAP7_75t_R register___U8226 ( .A(register__n3978), .Y(register__n4846) );
  INVx1_ASAP7_75t_R register___U8227 ( .A(register__n2847), .Y(register__n4847) );
  OA22x2_ASAP7_75t_R register___U8228 ( .A1(register__net64860), .A2(register__n1549), .B1(register__net104596), .B2(
        n1520), .Y(register__n12601) );
  OA22x2_ASAP7_75t_R register___U8229 ( .A1(register__n12194), .A2(register__n2851), .B1(register__n10022), .B2(register__n11750), 
        .Y(register__n13273) );
  INVx1_ASAP7_75t_R register___U8230 ( .A(register__n13273), .Y(register__n4853) );
  OA22x2_ASAP7_75t_R register___U8231 ( .A1(register__n12374), .A2(register__n104), .B1(register__n9915), .B2(register__n1618), 
        .Y(register__n12755) );
  INVx1_ASAP7_75t_R register___U8232 ( .A(register__n3607), .Y(register__n4854) );
  OA22x2_ASAP7_75t_R register___U8233 ( .A1(register__net64852), .A2(register__n665), .B1(register__net90077), .B2(
        n3746), .Y(register__n12826) );
  OA22x2_ASAP7_75t_R register___U8234 ( .A1(register__net63162), .A2(register__n2805), .B1(register__net97237), .B2(
        n4587), .Y(register__n12864) );
  INVx1_ASAP7_75t_R register___U8235 ( .A(register__n3396), .Y(register__n4855) );
  OA22x2_ASAP7_75t_R register___U8236 ( .A1(register__n12018), .A2(register__n3719), .B1(register__n10357), .B2(register__n1164), 
        .Y(register__n13385) );
  OA22x2_ASAP7_75t_R register___U8237 ( .A1(register__n12053), .A2(register__n576), .B1(register__n10456), .B2(register__n585), 
        .Y(register__n13230) );
  OA22x2_ASAP7_75t_R register___U8238 ( .A1(register__n12087), .A2(register__n1916), .B1(register__n10098), .B2(register__n11793), 
        .Y(register__n12909) );
  OA22x2_ASAP7_75t_R register___U8239 ( .A1(register__net64676), .A2(register__n956), .B1(register__n9728), .B2(register__n960), 
        .Y(register__n13031) );
  OA22x2_ASAP7_75t_R register___U8240 ( .A1(register__n3445), .A2(register__n11730), .B1(register__n9541), .B2(register__n1164), 
        .Y(register__n13375) );
  INVx1_ASAP7_75t_R register___U8241 ( .A(register__n3958), .Y(register__n4858) );
  OA22x2_ASAP7_75t_R register___U8242 ( .A1(register__n12117), .A2(register__n100), .B1(register__n9284), .B2(register__n11774), 
        .Y(register__n12967) );
  INVx1_ASAP7_75t_R register___U8243 ( .A(register__n12967), .Y(register__n4859) );
  OA22x2_ASAP7_75t_R register___U8244 ( .A1(register__net64000), .A2(register__n1755), .B1(register__net88584), .B2(
        n3821), .Y(register__n13132) );
  INVx1_ASAP7_75t_R register___U8245 ( .A(register__n3123), .Y(register__n4860) );
  OA22x2_ASAP7_75t_R register___U8246 ( .A1(register__net64014), .A2(register__n337), .B1(register__net96767), .B2(register__n68), 
        .Y(register__n12732) );
  OA22x2_ASAP7_75t_R register___U8247 ( .A1(register__net64006), .A2(register__n1416), .B1(register__net88412), .B2(
        n1419), .Y(register__n12995) );
  INVx1_ASAP7_75t_R register___U8248 ( .A(register__n3518), .Y(register__n4861) );
  BUFx2_ASAP7_75t_R register___U8249 ( .A(register__n10928), .Y(register__n4862) );
  BUFx2_ASAP7_75t_R register___U8250 ( .A(register__n8576), .Y(register__n4863) );
  INVx2_ASAP7_75t_R register___U8251 ( .A(register__n12331), .Y(register__n4864) );
  BUFx4f_ASAP7_75t_R register___U8252 ( .A(register__n12334), .Y(register__n12325) );
  BUFx12f_ASAP7_75t_R register___U8253 ( .A(register__n4834), .Y(register__n12331) );
  BUFx12f_ASAP7_75t_R register___U8254 ( .A(register__n3837), .Y(register__n4866) );
  BUFx4f_ASAP7_75t_R register___U8255 ( .A(register__n4195), .Y(register__n12037) );
  BUFx12f_ASAP7_75t_R register___U8256 ( .A(register__n4193), .Y(register__n12033) );
  BUFx2_ASAP7_75t_R register___U8257 ( .A(register__n4871), .Y(register__n4870) );
  BUFx2_ASAP7_75t_R register___U8258 ( .A(register__n13018), .Y(register__n4871) );
  INVx4_ASAP7_75t_R register___U8259 ( .A(register__n11865), .Y(register__n11864) );
  INVx5_ASAP7_75t_R register___U8260 ( .A(register__n11979), .Y(register__n11962) );
  BUFx2_ASAP7_75t_R register___U8261 ( .A(register__n4876), .Y(register__n4875) );
  BUFx2_ASAP7_75t_R register___U8262 ( .A(register__n12849), .Y(register__n4876) );
  BUFx2_ASAP7_75t_R register___U8263 ( .A(register__n4878), .Y(register__n4877) );
  BUFx2_ASAP7_75t_R register___U8264 ( .A(register__n4880), .Y(register__n4879) );
  BUFx2_ASAP7_75t_R register___U8265 ( .A(register__n13286), .Y(register__n4880) );
  BUFx2_ASAP7_75t_R register___U8266 ( .A(register__n4882), .Y(register__n4881) );
  BUFx2_ASAP7_75t_R register___U8267 ( .A(register__n13068), .Y(register__n4882) );
  BUFx2_ASAP7_75t_R register___U8268 ( .A(register__n13073), .Y(register__n4883) );
  BUFx2_ASAP7_75t_R register___U8269 ( .A(register__n4885), .Y(register__n4884) );
  BUFx2_ASAP7_75t_R register___U8270 ( .A(register__n4887), .Y(register__n4886) );
  BUFx2_ASAP7_75t_R register___U8271 ( .A(register__n4889), .Y(register__n4888) );
  BUFx2_ASAP7_75t_R register___U8272 ( .A(register__n13301), .Y(register__n4889) );
  BUFx2_ASAP7_75t_R register___U8273 ( .A(register__n4891), .Y(register__n4890) );
  BUFx2_ASAP7_75t_R register___U8274 ( .A(register__n4893), .Y(register__n4892) );
  BUFx2_ASAP7_75t_R register___U8275 ( .A(register__n13064), .Y(register__n4893) );
  INVx6_ASAP7_75t_R register___U8276 ( .A(register__n3678), .Y(register__n12170) );
  BUFx3_ASAP7_75t_R register___U8277 ( .A(register__n4895), .Y(register__n4894) );
  BUFx2_ASAP7_75t_R register___U8278 ( .A(register__n11528), .Y(register__n4895) );
  BUFx3_ASAP7_75t_R register___U8279 ( .A(register__n4897), .Y(register__n4896) );
  BUFx2_ASAP7_75t_R register___U8280 ( .A(register__n11529), .Y(register__n4897) );
  BUFx3_ASAP7_75t_R register___U8281 ( .A(register__n4899), .Y(register__n4898) );
  BUFx2_ASAP7_75t_R register___U8282 ( .A(register__n7297), .Y(register__n4900) );
  BUFx3_ASAP7_75t_R register___U8283 ( .A(register__n4902), .Y(register__n4901) );
  BUFx2_ASAP7_75t_R register___U8284 ( .A(register__n11184), .Y(register__n4902) );
  BUFx3_ASAP7_75t_R register___U8285 ( .A(register__n4904), .Y(register__n4903) );
  BUFx2_ASAP7_75t_R register___U8286 ( .A(register__n11185), .Y(register__n4904) );
  BUFx3_ASAP7_75t_R register___U8287 ( .A(register__n4906), .Y(register__n4905) );
  BUFx2_ASAP7_75t_R register___U8288 ( .A(register__n11118), .Y(register__n4906) );
  BUFx2_ASAP7_75t_R register___U8289 ( .A(register__n8264), .Y(register__n4909) );
  AO22x1_ASAP7_75t_R register___U8290 ( .A1(register__n9315), .A2(register__n3), .B1(register__n9417), .B2(register__n1579), .Y(
        n11120) );
  BUFx3_ASAP7_75t_R register___U8291 ( .A(register__n4915), .Y(register__n4914) );
  BUFx2_ASAP7_75t_R register___U8292 ( .A(register__n10623), .Y(register__n4915) );
  BUFx3_ASAP7_75t_R register___U8293 ( .A(register__n4917), .Y(register__n4916) );
  BUFx2_ASAP7_75t_R register___U8294 ( .A(register__n10624), .Y(register__n4917) );
  BUFx12f_ASAP7_75t_R register___U8295 ( .A(register__net64732), .Y(register__net64712) );
  BUFx12f_ASAP7_75t_R register___U8296 ( .A(register__n11808), .Y(register__n4920) );
  BUFx12f_ASAP7_75t_R register___U8297 ( .A(register__n3605), .Y(register__n11808) );
  BUFx2_ASAP7_75t_R register___U8298 ( .A(register__n10819), .Y(register__n4922) );
  BUFx3_ASAP7_75t_R register___U8299 ( .A(register__n4926), .Y(register__n4925) );
  BUFx2_ASAP7_75t_R register___U8300 ( .A(register__n10821), .Y(register__n4926) );
  BUFx2_ASAP7_75t_R register___U8301 ( .A(register__n7967), .Y(register__n4927) );
  BUFx3_ASAP7_75t_R register___U8302 ( .A(register__n4931), .Y(register__n4930) );
  BUFx2_ASAP7_75t_R register___U8303 ( .A(register__n10659), .Y(register__n4931) );
  BUFx3_ASAP7_75t_R register___U8304 ( .A(register__n4936), .Y(register__n4935) );
  BUFx2_ASAP7_75t_R register___U8305 ( .A(register__n10932), .Y(register__n4936) );
  BUFx3_ASAP7_75t_R register___U8306 ( .A(register__n10931), .Y(register__n4937) );
  BUFx3_ASAP7_75t_R register___U8307 ( .A(register__n4939), .Y(register__n4938) );
  BUFx2_ASAP7_75t_R register___U8308 ( .A(register__n10865), .Y(register__n4939) );
  BUFx3_ASAP7_75t_R register___U8309 ( .A(register__n4941), .Y(register__n4940) );
  BUFx2_ASAP7_75t_R register___U8310 ( .A(register__n10864), .Y(register__n4941) );
  BUFx3_ASAP7_75t_R register___U8311 ( .A(register__n4943), .Y(register__n4942) );
  BUFx3_ASAP7_75t_R register___U8312 ( .A(register__n4945), .Y(register__n4944) );
  BUFx2_ASAP7_75t_R register___U8313 ( .A(register__n10638), .Y(register__n4945) );
  BUFx2_ASAP7_75t_R register___U8314 ( .A(register__n28), .Y(register__n4946) );
  BUFx3_ASAP7_75t_R register___U8315 ( .A(register__n11057), .Y(register__n4949) );
  BUFx12f_ASAP7_75t_R register___U8316 ( .A(register__n5181), .Y(register__n11851) );
  BUFx3_ASAP7_75t_R register___U8317 ( .A(register__n6283), .Y(register__n4956) );
  BUFx2_ASAP7_75t_R register___U8318 ( .A(register__n9331), .Y(register__n4958) );
  BUFx2_ASAP7_75t_R register___U8319 ( .A(register__n9331), .Y(register__n4959) );
  BUFx3_ASAP7_75t_R register___U8320 ( .A(register__n10423), .Y(register__n4960) );
  BUFx4f_ASAP7_75t_R register___U8321 ( .A(register__n10423), .Y(register__n4961) );
  BUFx2_ASAP7_75t_R register___U8322 ( .A(register__n10423), .Y(register__n4962) );
  BUFx2_ASAP7_75t_R register___U8323 ( .A(register__n7685), .Y(register__n4963) );
  BUFx2_ASAP7_75t_R register___U8324 ( .A(register__n7687), .Y(register__n4965) );
  OR2x2_ASAP7_75t_R register___U8325 ( .A(register__n11846), .B(register__n11847), .Y(register__n7685) );
  BUFx12f_ASAP7_75t_R register___U8326 ( .A(register__n4838), .Y(register__n12244) );
  BUFx12f_ASAP7_75t_R register___U8327 ( .A(register__n4838), .Y(register__n12241) );
  BUFx3_ASAP7_75t_R register___U8328 ( .A(register__n4970), .Y(register__n4969) );
  BUFx2_ASAP7_75t_R register___U8329 ( .A(Reg_data[425]), .Y(register__n4970) );
  BUFx3_ASAP7_75t_R register___U8330 ( .A(register__net126193), .Y(register__net126192) );
  BUFx2_ASAP7_75t_R register___U8331 ( .A(Reg_data[746]), .Y(register__net126193) );
  BUFx3_ASAP7_75t_R register___U8332 ( .A(register__n4972), .Y(register__n4971) );
  BUFx2_ASAP7_75t_R register___U8333 ( .A(Reg_data[442]), .Y(register__n4972) );
  BUFx12f_ASAP7_75t_R register___U8334 ( .A(register__net139023), .Y(register__net63026) );
  BUFx12f_ASAP7_75t_R register___U8335 ( .A(register__net134980), .Y(register__net91923) );
  OA22x2_ASAP7_75t_R register___U8336 ( .A1(register__n12116), .A2(register__n955), .B1(register__n9879), .B2(register__n959), 
        .Y(register__n13026) );
  OA22x2_ASAP7_75t_R register___U8337 ( .A1(register__n99), .A2(register__n954), .B1(register__n9887), .B2(register__n958), .Y(
        n13022) );
  OA22x2_ASAP7_75t_R register___U8338 ( .A1(register__n12398), .A2(register__n1922), .B1(register__n6823), .B2(register__n1197), 
        .Y(register__n13091) );
  INVx1_ASAP7_75t_R register___U8339 ( .A(register__n3527), .Y(register__n4975) );
  INVx1_ASAP7_75t_R register___U8340 ( .A(register__n10744), .Y(register__n4976) );
  INVx1_ASAP7_75t_R register___U8341 ( .A(register__n3529), .Y(register__n4977) );
  INVx1_ASAP7_75t_R register___U8342 ( .A(register__n3108), .Y(register__n4978) );
  OA22x2_ASAP7_75t_R register___U8343 ( .A1(register__net62660), .A2(register__n954), .B1(register__n8125), .B2(register__n960), 
        .Y(register__n13010) );
  INVx1_ASAP7_75t_R register___U8344 ( .A(register__n3490), .Y(register__n4979) );
  OA22x2_ASAP7_75t_R register___U8345 ( .A1(register__n12052), .A2(register__n1049), .B1(register__n10024), .B2(register__n11745), 
        .Y(register__n13279) );
  INVx1_ASAP7_75t_R register___U8346 ( .A(register__n13279), .Y(register__n4980) );
  OA22x2_ASAP7_75t_R register___U8347 ( .A1(register__net64020), .A2(register__n119), .B1(register__net104592), .B2(
        n1527), .Y(register__n12593) );
  INVx1_ASAP7_75t_R register___U8348 ( .A(register__n3552), .Y(register__n4981) );
  OA22x2_ASAP7_75t_R register___U8349 ( .A1(register__n12346), .A2(register__n1793), .B1(register__n9917), .B2(register__n1620), 
        .Y(register__n12756) );
  OA22x2_ASAP7_75t_R register___U8350 ( .A1(register__net64936), .A2(register__n1069), .B1(register__n9947), .B2(register__n1992), 
        .Y(register__n12827) );
  OA22x2_ASAP7_75t_R register___U8351 ( .A1(register__n12257), .A2(register__n2806), .B1(register__n8708), .B2(register__n1936), 
        .Y(register__n12871) );
  INVx1_ASAP7_75t_R register___U8352 ( .A(register__n3484), .Y(register__n4982) );
  OA22x2_ASAP7_75t_R register___U8353 ( .A1(register__net64756), .A2(register__n1139), .B1(register__net97197), .B2(
        n1141), .Y(register__n13170) );
  INVx1_ASAP7_75t_R register___U8354 ( .A(register__n13170), .Y(register__n4983) );
  OA22x2_ASAP7_75t_R register___U8355 ( .A1(register__n12254), .A2(register__n577), .B1(register__n7337), .B2(register__n584), 
        .Y(register__n13220) );
  INVx1_ASAP7_75t_R register___U8356 ( .A(register__n3488), .Y(register__n4984) );
  OA22x2_ASAP7_75t_R register___U8357 ( .A1(register__n12143), .A2(register__n698), .B1(register__n10373), .B2(register__n669), 
        .Y(register__n13322) );
  OA22x2_ASAP7_75t_R register___U8358 ( .A1(register__net64344), .A2(register__n11881), .B1(register__net89613), .B2(
        n2843), .Y(register__n12907) );
  OA22x2_ASAP7_75t_R register___U8359 ( .A1(register__net64340), .A2(register__n954), .B1(register__net90661), .B2(register__n958), .Y(register__n13027) );
  OA22x2_ASAP7_75t_R register___U8360 ( .A1(register__n12086), .A2(register__n101), .B1(register__n9286), .B2(register__n11775), 
        .Y(register__n12970) );
  OA22x2_ASAP7_75t_R register___U8361 ( .A1(register__net63236), .A2(register__n11730), .B1(register__net88861), .B2(
        n1164), .Y(register__n13365) );
  INVx1_ASAP7_75t_R register___U8362 ( .A(register__n3369), .Y(register__n4987) );
  OA22x2_ASAP7_75t_R register___U8363 ( .A1(register__n12174), .A2(register__n337), .B1(register__n9794), .B2(register__n68), .Y(
        n12733) );
  OA22x2_ASAP7_75t_R register___U8364 ( .A1(register__n12420), .A2(register__n11730), .B1(register__n10391), .B2(register__n1164), 
        .Y(register__n13361) );
  INVx1_ASAP7_75t_R register___U8365 ( .A(register__n3971), .Y(register__n4988) );
  OA22x2_ASAP7_75t_R register___U8366 ( .A1(register__n12283), .A2(register__n1755), .B1(register__n8777), .B2(register__n3821), 
        .Y(register__n13128) );
  INVx1_ASAP7_75t_R register___U8367 ( .A(register__n3175), .Y(register__n4989) );
  INVx2_ASAP7_75t_R register___U8368 ( .A(register__n9549), .Y(register__n10743) );
  BUFx3_ASAP7_75t_R register___U8369 ( .A(register__n4992), .Y(register__n4991) );
  BUFx2_ASAP7_75t_R register___U8370 ( .A(register__n10677), .Y(register__n4992) );
  BUFx2_ASAP7_75t_R register___U8371 ( .A(register__n10944), .Y(register__n4993) );
  BUFx2_ASAP7_75t_R register___U8372 ( .A(register__n6828), .Y(register__n4996) );
  BUFx12f_ASAP7_75t_R register___U8373 ( .A(register__n5345), .Y(register__n12355) );
  BUFx2_ASAP7_75t_R register___U8374 ( .A(register__n5003), .Y(register__n5002) );
  BUFx2_ASAP7_75t_R register___U8375 ( .A(register__n12671), .Y(register__n5003) );
  BUFx2_ASAP7_75t_R register___U8376 ( .A(register__n5005), .Y(register__n5004) );
  BUFx2_ASAP7_75t_R register___U8377 ( .A(register__n5012), .Y(register__n5011) );
  BUFx2_ASAP7_75t_R register___U8378 ( .A(register__n10546), .Y(register__n5015) );
  BUFx2_ASAP7_75t_R register___U8379 ( .A(register__n8566), .Y(register__n5016) );
  BUFx3_ASAP7_75t_R register___U8380 ( .A(register__n5018), .Y(register__n5017) );
  BUFx2_ASAP7_75t_R register___U8381 ( .A(register__n10543), .Y(register__n5018) );
  BUFx3_ASAP7_75t_R register___U8382 ( .A(register__n5020), .Y(register__n5019) );
  BUFx2_ASAP7_75t_R register___U8383 ( .A(register__n10545), .Y(register__n5020) );
  BUFx3_ASAP7_75t_R register___U8384 ( .A(register__n10946), .Y(register__n5021) );
  BUFx3_ASAP7_75t_R register___U8385 ( .A(register__n10948), .Y(register__n5022) );
  BUFx3_ASAP7_75t_R register___U8386 ( .A(register__n11145), .Y(register__n5025) );
  AO22x1_ASAP7_75t_R register___U8387 ( .A1(register__n8126), .A2(register__n1909), .B1(register__n10467), .B2(register__n381), 
        .Y(register__n11147) );
  BUFx3_ASAP7_75t_R register___U8388 ( .A(register__n5029), .Y(register__n5028) );
  BUFx2_ASAP7_75t_R register___U8389 ( .A(register__n10751), .Y(register__n5029) );
  BUFx3_ASAP7_75t_R register___U8390 ( .A(register__n5307), .Y(register__n8635) );
  BUFx3_ASAP7_75t_R register___U8391 ( .A(register__n5033), .Y(register__n5032) );
  BUFx2_ASAP7_75t_R register___U8392 ( .A(register__n11030), .Y(register__n5033) );
  BUFx12f_ASAP7_75t_R register___U8393 ( .A(register__net140271), .Y(register__net64384) );
  BUFx12f_ASAP7_75t_R register___U8394 ( .A(register__n12240), .Y(register__n12242) );
  BUFx12f_ASAP7_75t_R register___U8395 ( .A(register__n4837), .Y(register__n12240) );
  BUFx3_ASAP7_75t_R register___U8396 ( .A(register__n5037), .Y(register__n5036) );
  BUFx2_ASAP7_75t_R register___U8397 ( .A(register__n11265), .Y(register__n5037) );
  INVx2_ASAP7_75t_R register___U8398 ( .A(register__n7668), .Y(register__n5038) );
  BUFx3_ASAP7_75t_R register___U8399 ( .A(register__n5040), .Y(register__n5039) );
  BUFx2_ASAP7_75t_R register___U8400 ( .A(register__n11264), .Y(register__n5040) );
  BUFx12f_ASAP7_75t_R register___U8401 ( .A(register__n8246), .Y(register__n5042) );
  BUFx12f_ASAP7_75t_R register___U8402 ( .A(register__n5525), .Y(register__n11835) );
  BUFx3_ASAP7_75t_R register___U8403 ( .A(register__n7389), .Y(register__n5046) );
  BUFx12f_ASAP7_75t_R register___U8404 ( .A(register__n11875), .Y(register__n11874) );
  BUFx6f_ASAP7_75t_R register___U8405 ( .A(register__n4194), .Y(register__n12042) );
  BUFx4f_ASAP7_75t_R register___U8406 ( .A(register__n3992), .Y(register__n12046) );
  BUFx4f_ASAP7_75t_R register___U8407 ( .A(register__n3992), .Y(register__n12047) );
  INVx2_ASAP7_75t_R register___U8408 ( .A(register__net63016), .Y(register__net62996) );
  BUFx12f_ASAP7_75t_R register___U8409 ( .A(register__net129690), .Y(register__net63046) );
  OA22x2_ASAP7_75t_R register___U8410 ( .A1(register__n12463), .A2(register__n117), .B1(register__n10389), .B2(register__n1663), 
        .Y(register__n12636) );
  OA22x2_ASAP7_75t_R register___U8411 ( .A1(register__net64836), .A2(register__n11868), .B1(register__net89861), .B2(
        n11751), .Y(register__n13280) );
  OA22x2_ASAP7_75t_R register___U8412 ( .A1(register__n12291), .A2(register__n3022), .B1(register__n7132), .B2(register__n1600), 
        .Y(register__n12700) );
  OA22x2_ASAP7_75t_R register___U8413 ( .A1(register__n12371), .A2(register__n462), .B1(register__n9987), .B2(register__n467), 
        .Y(register__n12927) );
  INVx1_ASAP7_75t_R register___U8414 ( .A(register__n3684), .Y(register__n5052) );
  OA22x2_ASAP7_75t_R register___U8415 ( .A1(register__net64840), .A2(register__n103), .B1(register__net97193), .B2(
        n1149), .Y(register__n13171) );
  OA22x2_ASAP7_75t_R register___U8416 ( .A1(register__net64754), .A2(register__n577), .B1(register__net89777), .B2(register__n581), .Y(register__n13232) );
  OA22x2_ASAP7_75t_R register___U8417 ( .A1(register__net64762), .A2(register__n101), .B1(register__net93741), .B2(
        n11777), .Y(register__n12973) );
  INVx1_ASAP7_75t_R register___U8418 ( .A(register__n12973), .Y(register__n5053) );
  OA22x2_ASAP7_75t_R register___U8419 ( .A1(register__net63322), .A2(register__n698), .B1(register__n9551), .B2(register__n679), 
        .Y(register__n13314) );
  OA22x2_ASAP7_75t_R register___U8420 ( .A1(register__net64684), .A2(register__n1069), .B1(register__n10185), .B2(register__n81), 
        .Y(register__n12824) );
  INVx1_ASAP7_75t_R register___U8421 ( .A(register__n3520), .Y(register__n5054) );
  OA22x2_ASAP7_75t_R register___U8422 ( .A1(register__net64420), .A2(register__n339), .B1(register__net96863), .B2(register__n343), .Y(register__n12737) );
  INVx1_ASAP7_75t_R register___U8423 ( .A(register__n3775), .Y(register__n5055) );
  OA22x2_ASAP7_75t_R register___U8424 ( .A1(register__net64420), .A2(register__n11730), .B1(register__net88821), .B2(
        n1164), .Y(register__n13379) );
  INVx1_ASAP7_75t_R register___U8425 ( .A(register__n3402), .Y(register__n5056) );
  OA22x2_ASAP7_75t_R register___U8426 ( .A1(register__net64424), .A2(register__n952), .B1(register__net88404), .B2(register__n959), .Y(register__n13028) );
  OA22x2_ASAP7_75t_R register___U8427 ( .A1(register__net63328), .A2(register__n1755), .B1(register__n9843), .B2(register__n3821), 
        .Y(register__n13124) );
  INVx1_ASAP7_75t_R register___U8428 ( .A(register__n3226), .Y(register__n5057) );
  OA22x2_ASAP7_75t_R register___U8429 ( .A1(register__net143255), .A2(register__n1415), .B1(register__n9845), .B2(register__n1419), .Y(register__n12987) );
  INVx1_ASAP7_75t_R register___U8430 ( .A(register__n3556), .Y(register__n5058) );
  INVx2_ASAP7_75t_R register___U8431 ( .A(register__n9545), .Y(register__n11587) );
  BUFx3_ASAP7_75t_R register___U8432 ( .A(register__n5060), .Y(register__n5059) );
  BUFx2_ASAP7_75t_R register___U8433 ( .A(register__n11254), .Y(register__n5060) );
  BUFx2_ASAP7_75t_R register___U8434 ( .A(register__n8234), .Y(register__n5061) );
  AO22x1_ASAP7_75t_R register___U8435 ( .A1(register__net90925), .A2(register__n3), .B1(register__net90017), .B2(register__n1578), 
        .Y(register__n11012) );
  BUFx3_ASAP7_75t_R register___U8436 ( .A(register__n5063), .Y(register__n5062) );
  BUFx2_ASAP7_75t_R register___U8437 ( .A(register__n10949), .Y(register__n5063) );
  BUFx3_ASAP7_75t_R register___U8438 ( .A(register__n5065), .Y(register__n5064) );
  BUFx2_ASAP7_75t_R register___U8439 ( .A(register__n10582), .Y(register__n5065) );
  BUFx3_ASAP7_75t_R register___U8440 ( .A(register__n5067), .Y(register__n5066) );
  BUFx2_ASAP7_75t_R register___U8441 ( .A(register__n10778), .Y(register__n5067) );
  BUFx3_ASAP7_75t_R register___U8442 ( .A(register__n5071), .Y(register__n5070) );
  BUFx2_ASAP7_75t_R register___U8443 ( .A(register__n10649), .Y(register__n5071) );
  BUFx3_ASAP7_75t_R register___U8444 ( .A(register__n5073), .Y(register__n5072) );
  BUFx2_ASAP7_75t_R register___U8445 ( .A(register__n11652), .Y(register__n5073) );
  BUFx2_ASAP7_75t_R register___U8446 ( .A(register__n5076), .Y(register__n5075) );
  BUFx2_ASAP7_75t_R register___U8447 ( .A(register__n12757), .Y(register__n5076) );
  BUFx2_ASAP7_75t_R register___U8448 ( .A(register__n5078), .Y(register__n5077) );
  BUFx2_ASAP7_75t_R register___U8449 ( .A(register__n13045), .Y(register__n5078) );
  BUFx2_ASAP7_75t_R register___U8450 ( .A(register__n5084), .Y(register__n5083) );
  BUFx2_ASAP7_75t_R register___U8451 ( .A(register__n13060), .Y(register__n5084) );
  BUFx2_ASAP7_75t_R register___U8452 ( .A(register__n5086), .Y(register__n5085) );
  BUFx2_ASAP7_75t_R register___U8453 ( .A(register__n13056), .Y(register__n5086) );
  BUFx2_ASAP7_75t_R register___U8454 ( .A(register__n5090), .Y(register__n5089) );
  BUFx2_ASAP7_75t_R register___U8455 ( .A(register__n12654), .Y(register__n5090) );
  BUFx2_ASAP7_75t_R register___U8456 ( .A(register__n12653), .Y(register__n5092) );
  BUFx2_ASAP7_75t_R register___U8457 ( .A(register__n5096), .Y(register__n5095) );
  BUFx2_ASAP7_75t_R register___U8458 ( .A(register__n12751), .Y(register__n5096) );
  BUFx2_ASAP7_75t_R register___U8459 ( .A(register__n5098), .Y(register__n5097) );
  BUFx2_ASAP7_75t_R register___U8460 ( .A(register__n5100), .Y(register__n5099) );
  BUFx2_ASAP7_75t_R register___U8461 ( .A(register__n12649), .Y(register__n5100) );
  BUFx3_ASAP7_75t_R register___U8462 ( .A(register__n5105), .Y(register__n5104) );
  BUFx2_ASAP7_75t_R register___U8463 ( .A(register__n10653), .Y(register__n5105) );
  BUFx2_ASAP7_75t_R register___U8464 ( .A(register__n10654), .Y(register__n5106) );
  BUFx2_ASAP7_75t_R register___U8465 ( .A(register__n7004), .Y(register__n5107) );
  BUFx3_ASAP7_75t_R register___U8466 ( .A(register__n5111), .Y(register__n5110) );
  BUFx2_ASAP7_75t_R register___U8467 ( .A(register__n11364), .Y(register__n5111) );
  BUFx3_ASAP7_75t_R register___U8468 ( .A(register__n5113), .Y(register__n5112) );
  BUFx2_ASAP7_75t_R register___U8469 ( .A(register__n11613), .Y(register__n5113) );
  BUFx3_ASAP7_75t_R register___U8470 ( .A(register__n5115), .Y(register__n5114) );
  BUFx2_ASAP7_75t_R register___U8471 ( .A(register__n11616), .Y(register__n5115) );
  BUFx12f_ASAP7_75t_R register___U8472 ( .A(register__n3846), .Y(register__n12012) );
  BUFx2_ASAP7_75t_R register___U8473 ( .A(register__n8328), .Y(register__n5117) );
  BUFx2_ASAP7_75t_R register___U8474 ( .A(register__n8329), .Y(register__n5118) );
  BUFx12f_ASAP7_75t_R register___U8475 ( .A(register__net64360), .Y(register__net64382) );
  BUFx3_ASAP7_75t_R register___U8476 ( .A(register__n5120), .Y(register__n5119) );
  BUFx3_ASAP7_75t_R register___U8477 ( .A(register__n5122), .Y(register__n5121) );
  BUFx2_ASAP7_75t_R register___U8478 ( .A(register__n11432), .Y(register__n5122) );
  BUFx3_ASAP7_75t_R register___U8479 ( .A(register__n11431), .Y(register__n5123) );
  BUFx4f_ASAP7_75t_R register___U8480 ( .A(register__n5123), .Y(register__n7674) );
  BUFx3_ASAP7_75t_R register___U8481 ( .A(register__n5127), .Y(register__n5126) );
  BUFx2_ASAP7_75t_R register___U8482 ( .A(register__n10527), .Y(register__n5127) );
  BUFx2_ASAP7_75t_R register___U8483 ( .A(register__n8305), .Y(register__n5129) );
  BUFx3_ASAP7_75t_R register___U8484 ( .A(register__n5131), .Y(register__n5130) );
  BUFx2_ASAP7_75t_R register___U8485 ( .A(register__n11000), .Y(register__n5131) );
  BUFx3_ASAP7_75t_R register___U8486 ( .A(register__n5133), .Y(register__n5132) );
  BUFx2_ASAP7_75t_R register___U8487 ( .A(register__n10999), .Y(register__n5133) );
  BUFx3_ASAP7_75t_R register___U8488 ( .A(register__n5135), .Y(register__n5134) );
  BUFx2_ASAP7_75t_R register___U8489 ( .A(register__n10912), .Y(register__n5135) );
  BUFx3_ASAP7_75t_R register___U8490 ( .A(register__n5137), .Y(register__n5136) );
  BUFx2_ASAP7_75t_R register___U8491 ( .A(register__n10911), .Y(register__n5137) );
  BUFx3_ASAP7_75t_R register___U8492 ( .A(register__n5139), .Y(register__n5138) );
  BUFx2_ASAP7_75t_R register___U8493 ( .A(register__n10758), .Y(register__n5139) );
  BUFx3_ASAP7_75t_R register___U8494 ( .A(register__n5141), .Y(register__n5140) );
  BUFx2_ASAP7_75t_R register___U8495 ( .A(register__n10703), .Y(register__n5141) );
  BUFx3_ASAP7_75t_R register___U8496 ( .A(register__n5143), .Y(register__n5142) );
  BUFx2_ASAP7_75t_R register___U8497 ( .A(register__n10702), .Y(register__n5143) );
  BUFx2_ASAP7_75t_R register___U8498 ( .A(register__n9), .Y(register__n5144) );
  BUFx3_ASAP7_75t_R register___U8499 ( .A(register__n5146), .Y(register__n5145) );
  BUFx2_ASAP7_75t_R register___U8500 ( .A(register__n10844), .Y(register__n5146) );
  BUFx3_ASAP7_75t_R register___U8501 ( .A(register__n5148), .Y(register__n5147) );
  BUFx2_ASAP7_75t_R register___U8502 ( .A(register__n10843), .Y(register__n5148) );
  BUFx3_ASAP7_75t_R register___U8503 ( .A(register__n11303), .Y(register__n5149) );
  INVx2_ASAP7_75t_R register___U8504 ( .A(register__n70), .Y(register__n5150) );
  BUFx3_ASAP7_75t_R register___U8505 ( .A(register__n5152), .Y(register__n5151) );
  BUFx3_ASAP7_75t_R register___U8506 ( .A(register__n5154), .Y(register__n5153) );
  BUFx2_ASAP7_75t_R register___U8507 ( .A(register__n11124), .Y(register__n5154) );
  BUFx3_ASAP7_75t_R register___U8508 ( .A(register__n5156), .Y(register__n5155) );
  BUFx3_ASAP7_75t_R register___U8509 ( .A(register__n5159), .Y(register__n5158) );
  BUFx2_ASAP7_75t_R register___U8510 ( .A(register__n10805), .Y(register__n5159) );
  BUFx2_ASAP7_75t_R register___U8511 ( .A(register__n8312), .Y(register__n5161) );
  BUFx3_ASAP7_75t_R register___U8512 ( .A(register__n10804), .Y(register__n5162) );
  BUFx3_ASAP7_75t_R register___U8513 ( .A(register__n5164), .Y(register__n5163) );
  BUFx2_ASAP7_75t_R register___U8514 ( .A(register__n11016), .Y(register__n5164) );
  BUFx3_ASAP7_75t_R register___U8515 ( .A(register__n5166), .Y(register__n5165) );
  BUFx2_ASAP7_75t_R register___U8516 ( .A(register__n11015), .Y(register__n5166) );
  BUFx2_ASAP7_75t_R register___U8517 ( .A(register__n8325), .Y(register__n5169) );
  BUFx12f_ASAP7_75t_R register___U8518 ( .A(register__n5172), .Y(register__n5171) );
  BUFx3_ASAP7_75t_R register___U8519 ( .A(register__n9591), .Y(register__n5174) );
  BUFx4f_ASAP7_75t_R register___U8520 ( .A(register__n9591), .Y(register__n5175) );
  BUFx3_ASAP7_75t_R register___U8521 ( .A(register__net105810), .Y(register__net123812) );
  BUFx3_ASAP7_75t_R register___U8522 ( .A(register__n8485), .Y(register__n5176) );
  BUFx3_ASAP7_75t_R register___U8523 ( .A(register__n7534), .Y(register__n5177) );
  BUFx3_ASAP7_75t_R register___U8524 ( .A(register__n8183), .Y(register__n5178) );
  BUFx3_ASAP7_75t_R register___U8525 ( .A(register__n7853), .Y(register__n5179) );
  BUFx12f_ASAP7_75t_R register___U8526 ( .A(register__n10334), .Y(register__n5180) );
  OR2x2_ASAP7_75t_R register___U8527 ( .A(register__n1422), .B(register__n4963), .Y(register__n7686) );
  OR2x2_ASAP7_75t_R register___U8528 ( .A(register__n1489), .B(register__n1282), .Y(register__n7687) );
  AND3x1_ASAP7_75t_R register___U8529 ( .A(register__n4376), .B(register__n12518), .C(register__n12519), .Y(register__n12517) );
  INVx6_ASAP7_75t_R register___U8530 ( .A(register__n781), .Y(register__n5185) );
  BUFx12f_ASAP7_75t_R register___U8531 ( .A(register__n5185), .Y(register__n12246) );
  BUFx3_ASAP7_75t_R register___U8532 ( .A(register__n5187), .Y(register__n5186) );
  BUFx2_ASAP7_75t_R register___U8533 ( .A(Reg_data[950]), .Y(register__n5187) );
  BUFx3_ASAP7_75t_R register___U8534 ( .A(register__n5189), .Y(register__n5188) );
  BUFx2_ASAP7_75t_R register___U8535 ( .A(Reg_data[948]), .Y(register__n5189) );
  BUFx2_ASAP7_75t_R register___U8536 ( .A(register__n9583), .Y(register__n5190) );
  BUFx3_ASAP7_75t_R register___U8537 ( .A(register__n9583), .Y(register__n5191) );
  BUFx4f_ASAP7_75t_R register___U8538 ( .A(register__n9583), .Y(register__n5192) );
  BUFx3_ASAP7_75t_R register___U8539 ( .A(register__n5194), .Y(register__n5193) );
  BUFx2_ASAP7_75t_R register___U8540 ( .A(Reg_data[944]), .Y(register__n5194) );
  BUFx3_ASAP7_75t_R register___U8541 ( .A(register__net123676), .Y(register__net123675) );
  BUFx2_ASAP7_75t_R register___U8542 ( .A(Reg_data[933]), .Y(register__net123676) );
  BUFx3_ASAP7_75t_R register___U8543 ( .A(register__n5196), .Y(register__n5195) );
  BUFx2_ASAP7_75t_R register___U8544 ( .A(Reg_data[929]), .Y(register__n5196) );
  BUFx3_ASAP7_75t_R register___U8545 ( .A(register__n8341), .Y(register__n5197) );
  BUFx4f_ASAP7_75t_R register___U8546 ( .A(register__n8341), .Y(register__n5198) );
  BUFx2_ASAP7_75t_R register___U8547 ( .A(register__n8341), .Y(register__n5199) );
  BUFx3_ASAP7_75t_R register___U8548 ( .A(register__n5201), .Y(register__n5200) );
  BUFx2_ASAP7_75t_R register___U8549 ( .A(Reg_data[725]), .Y(register__n5201) );
  BUFx3_ASAP7_75t_R register___U8550 ( .A(register__n5203), .Y(register__n5202) );
  BUFx2_ASAP7_75t_R register___U8551 ( .A(Reg_data[712]), .Y(register__n5203) );
  BUFx3_ASAP7_75t_R register___U8552 ( .A(register__n5205), .Y(register__n5204) );
  BUFx2_ASAP7_75t_R register___U8553 ( .A(Reg_data[178]), .Y(register__n5205) );
  BUFx3_ASAP7_75t_R register___U8554 ( .A(register__n10004), .Y(register__n5206) );
  BUFx4f_ASAP7_75t_R register___U8555 ( .A(register__n10004), .Y(register__n5207) );
  BUFx2_ASAP7_75t_R register___U8556 ( .A(register__n10004), .Y(register__n5208) );
  BUFx3_ASAP7_75t_R register___U8557 ( .A(register__n5210), .Y(register__n5209) );
  BUFx2_ASAP7_75t_R register___U8558 ( .A(Reg_data[942]), .Y(register__n5210) );
  BUFx2_ASAP7_75t_R register___U8559 ( .A(register__n9806), .Y(register__n5211) );
  BUFx3_ASAP7_75t_R register___U8560 ( .A(register__n9806), .Y(register__n5212) );
  BUFx4f_ASAP7_75t_R register___U8561 ( .A(register__n3251), .Y(register__n5214) );
  BUFx2_ASAP7_75t_R register___U8562 ( .A(Reg_data[187]), .Y(register__n5215) );
  BUFx6f_ASAP7_75t_R register___U8563 ( .A(register__n5214), .Y(register__n10267) );
  INVx2_ASAP7_75t_R register___U8564 ( .A(register__n12035), .Y(register__n12019) );
  BUFx4f_ASAP7_75t_R register___U8565 ( .A(register__n4866), .Y(register__n12035) );
  BUFx12f_ASAP7_75t_R register___U8566 ( .A(register__net105198), .Y(register__net123601) );
  OA22x2_ASAP7_75t_R register___U8567 ( .A1(register__n12235), .A2(register__n1657), .B1(register__n9517), .B2(register__n1670), 
        .Y(register__n12646) );
  INVx1_ASAP7_75t_R register___U8568 ( .A(register__n4403), .Y(register__n5216) );
  OA22x2_ASAP7_75t_R register___U8569 ( .A1(register__net62842), .A2(register__n116), .B1(register__net88752), .B2(
        n1679), .Y(register__n12637) );
  OA22x2_ASAP7_75t_R register___U8570 ( .A1(register__net62660), .A2(register__n890), .B1(register__n6923), .B2(register__n898), 
        .Y(register__n13038) );
  OA22x2_ASAP7_75t_R register___U8571 ( .A1(register__net64416), .A2(register__n1793), .B1(register__net115978), .B2(
        n1623), .Y(register__n12766) );
  INVx1_ASAP7_75t_R register___U8572 ( .A(register__n3779), .Y(register__n5220) );
  OA22x2_ASAP7_75t_R register___U8573 ( .A1(register__n12290), .A2(register__n1792), .B1(register__n6950), .B2(register__n1642), 
        .Y(register__n12758) );
  INVx1_ASAP7_75t_R register___U8574 ( .A(register__n12758), .Y(register__n5221) );
  OA22x2_ASAP7_75t_R register___U8575 ( .A1(register__net62838), .A2(register__n1643), .B1(register__net94787), .B2(
        n1634), .Y(register__n12748) );
  INVx1_ASAP7_75t_R register___U8576 ( .A(register__n4539), .Y(register__n5222) );
  BUFx12f_ASAP7_75t_R register___U8577 ( .A(register__n3841), .Y(register__n5225) );
  BUFx12f_ASAP7_75t_R register___U8578 ( .A(register__n5224), .Y(register__n12470) );
  BUFx4f_ASAP7_75t_R register___U8579 ( .A(register__n3215), .Y(register__n12467) );
  INVx1_ASAP7_75t_R register___U8580 ( .A(register__n3137), .Y(register__n5228) );
  INVx1_ASAP7_75t_R register___U8581 ( .A(register__n3139), .Y(register__n5229) );
  INVx1_ASAP7_75t_R register___U8582 ( .A(register__n4115), .Y(register__n5231) );
  OA22x2_ASAP7_75t_R register___U8583 ( .A1(register__n11951), .A2(register__n2851), .B1(register__n8349), .B2(register__n3438), 
        .Y(register__n13284) );
  OA22x2_ASAP7_75t_R register___U8584 ( .A1(register__n12203), .A2(register__n3022), .B1(register__n7328), .B2(register__n1586), 
        .Y(register__n12703) );
  OA22x2_ASAP7_75t_R register___U8585 ( .A1(register__n11960), .A2(register__n1792), .B1(register__n9325), .B2(register__n1631), 
        .Y(register__n12775) );
  INVx1_ASAP7_75t_R register___U8586 ( .A(register__n4499), .Y(register__n5235) );
  OA22x2_ASAP7_75t_R register___U8587 ( .A1(register__net64850), .A2(register__n2821), .B1(register__net97225), .B2(
        n1932), .Y(register__n12882) );
  OA22x2_ASAP7_75t_R register___U8588 ( .A1(register__n12340), .A2(register__n461), .B1(register__n9989), .B2(register__n463), 
        .Y(register__n12928) );
  OA22x2_ASAP7_75t_R register___U8589 ( .A1(register__n11953), .A2(register__n1137), .B1(register__n7986), .B2(register__n1150), 
        .Y(register__n13175) );
  OA22x2_ASAP7_75t_R register___U8590 ( .A1(register__net64838), .A2(register__n578), .B1(register__net89773), .B2(register__n589), .Y(register__n13233) );
  OA22x2_ASAP7_75t_R register___U8591 ( .A1(register__net64920), .A2(register__n101), .B1(register__n9290), .B2(register__n10517), 
        .Y(register__n12975) );
  INVx1_ASAP7_75t_R register___U8592 ( .A(register__n3083), .Y(register__n5238) );
  OA22x2_ASAP7_75t_R register___U8593 ( .A1(register__net63994), .A2(register__n700), .B1(register__net88857), .B2(register__n677), .Y(register__n13321) );
  OA22x2_ASAP7_75t_R register___U8594 ( .A1(register__net63000), .A2(register__n1974), .B1(register__n10426), .B2(
        n11883), .Y(register__n12892) );
  INVx1_ASAP7_75t_R register___U8595 ( .A(register__n3048), .Y(register__n5239) );
  OA22x2_ASAP7_75t_R register___U8596 ( .A1(register__n12173), .A2(register__n665), .B1(register__n10214), .B2(register__n81), 
        .Y(register__n12817) );
  INVx1_ASAP7_75t_R register___U8597 ( .A(register__n3773), .Y(register__n5240) );
  OA22x2_ASAP7_75t_R register___U8598 ( .A1(register__n12121), .A2(register__n337), .B1(register__n8775), .B2(register__n346), 
        .Y(register__n12735) );
  OA22x2_ASAP7_75t_R register___U8599 ( .A1(register__net63320), .A2(register__n11730), .B1(register__n10399), .B2(
        n1164), .Y(register__n13366) );
  INVx1_ASAP7_75t_R register___U8600 ( .A(register__n3434), .Y(register__n5242) );
  OA22x2_ASAP7_75t_R register___U8601 ( .A1(register__n2132), .A2(register__n1755), .B1(register__n9847), .B2(register__n3334), 
        .Y(register__n13138) );
  OA22x2_ASAP7_75t_R register___U8602 ( .A1(register__n12399), .A2(register__n954), .B1(register__n9871), .B2(register__n959), 
        .Y(register__n13014) );
  INVx1_ASAP7_75t_R register___U8603 ( .A(register__n3558), .Y(register__n5243) );
  OA22x2_ASAP7_75t_R register___U8604 ( .A1(register__n12400), .A2(register__n1416), .B1(register__n9873), .B2(register__n1418), 
        .Y(register__n12984) );
  INVx1_ASAP7_75t_R register___U8605 ( .A(register__n4090), .Y(register__n5244) );
  INVx2_ASAP7_75t_R register___U8606 ( .A(register__n9441), .Y(register__n10600) );
  INVx2_ASAP7_75t_R register___U8607 ( .A(register__n10339), .Y(register__n11180) );
  INVx2_ASAP7_75t_R register___U8608 ( .A(register__n7997), .Y(register__n11352) );
  BUFx2_ASAP7_75t_R register___U8609 ( .A(register__n10981), .Y(register__n5246) );
  BUFx4f_ASAP7_75t_R register___U8610 ( .A(register__n9161), .Y(register__n6780) );
  BUFx3_ASAP7_75t_R register___U8611 ( .A(register__n5249), .Y(register__n5248) );
  BUFx2_ASAP7_75t_R register___U8612 ( .A(register__n11190), .Y(register__n5249) );
  BUFx3_ASAP7_75t_R register___U8613 ( .A(register__n5251), .Y(register__n5250) );
  BUFx2_ASAP7_75t_R register___U8614 ( .A(register__n11168), .Y(register__n5251) );
  BUFx2_ASAP7_75t_R register___U8615 ( .A(register__n5664), .Y(register__n5252) );
  BUFx3_ASAP7_75t_R register___U8616 ( .A(register__n5254), .Y(register__n5253) );
  BUFx2_ASAP7_75t_R register___U8617 ( .A(register__n10972), .Y(register__n5254) );
  BUFx3_ASAP7_75t_R register___U8618 ( .A(register__n5257), .Y(register__n5256) );
  BUFx2_ASAP7_75t_R register___U8619 ( .A(register__n11400), .Y(register__n5257) );
  BUFx2_ASAP7_75t_R register___U8620 ( .A(register__n8569), .Y(register__n5260) );
  BUFx3_ASAP7_75t_R register___U8621 ( .A(register__n5262), .Y(register__n5261) );
  BUFx2_ASAP7_75t_R register___U8622 ( .A(register__n10993), .Y(register__n5262) );
  BUFx2_ASAP7_75t_R register___U8623 ( .A(register__n8570), .Y(register__n5263) );
  AO22x1_ASAP7_75t_R register___U8624 ( .A1(register__n9764), .A2(register__n155), .B1(register__n10257), .B2(register__n381), 
        .Y(register__n10993) );
  BUFx3_ASAP7_75t_R register___U8625 ( .A(register__n5267), .Y(register__n5266) );
  BUFx2_ASAP7_75t_R register___U8626 ( .A(register__n11594), .Y(register__n5267) );
  BUFx2_ASAP7_75t_R register___U8627 ( .A(register__n5269), .Y(register__n5268) );
  BUFx6f_ASAP7_75t_R register___U8628 ( .A(register__n3469), .Y(register__n12207) );
  BUFx3_ASAP7_75t_R register___U8629 ( .A(register__n5275), .Y(register__n5274) );
  BUFx2_ASAP7_75t_R register___U8630 ( .A(register__n10675), .Y(register__n5275) );
  BUFx2_ASAP7_75t_R register___U8631 ( .A(register__n10674), .Y(register__n5278) );
  BUFx3_ASAP7_75t_R register___U8632 ( .A(register__n5280), .Y(register__n5279) );
  BUFx2_ASAP7_75t_R register___U8633 ( .A(register__n10632), .Y(register__n5280) );
  BUFx2_ASAP7_75t_R register___U8634 ( .A(register__n6417), .Y(register__n5281) );
  BUFx3_ASAP7_75t_R register___U8635 ( .A(register__n5283), .Y(register__n5282) );
  BUFx2_ASAP7_75t_R register___U8636 ( .A(register__n10631), .Y(register__n5283) );
  BUFx3_ASAP7_75t_R register___U8637 ( .A(register__n5285), .Y(register__n5284) );
  BUFx2_ASAP7_75t_R register___U8638 ( .A(register__n10729), .Y(register__n5285) );
  BUFx3_ASAP7_75t_R register___U8639 ( .A(register__n5287), .Y(register__n5286) );
  BUFx2_ASAP7_75t_R register___U8640 ( .A(register__n10856), .Y(register__n5287) );
  BUFx3_ASAP7_75t_R register___U8641 ( .A(register__n5291), .Y(register__n5290) );
  BUFx2_ASAP7_75t_R register___U8642 ( .A(register__n11074), .Y(register__n5291) );
  BUFx3_ASAP7_75t_R register___U8643 ( .A(register__n5293), .Y(register__n5292) );
  BUFx2_ASAP7_75t_R register___U8644 ( .A(register__n11075), .Y(register__n5293) );
  BUFx3_ASAP7_75t_R register___U8645 ( .A(register__n5295), .Y(register__n5294) );
  BUFx2_ASAP7_75t_R register___U8646 ( .A(register__n11076), .Y(register__n5295) );
  BUFx3_ASAP7_75t_R register___U8647 ( .A(register__n5297), .Y(register__n5296) );
  BUFx2_ASAP7_75t_R register___U8648 ( .A(register__n11093), .Y(register__n5297) );
  BUFx2_ASAP7_75t_R register___U8649 ( .A(register__n11094), .Y(register__n5298) );
  BUFx3_ASAP7_75t_R register___U8650 ( .A(register__n5300), .Y(register__n5299) );
  BUFx2_ASAP7_75t_R register___U8651 ( .A(register__n11095), .Y(register__n5300) );
  BUFx3_ASAP7_75t_R register___U8652 ( .A(register__n5303), .Y(register__n5302) );
  BUFx2_ASAP7_75t_R register___U8653 ( .A(register__n11690), .Y(register__n5303) );
  INVx1_ASAP7_75t_R register___U8654 ( .A(register__n8635), .Y(register__n5304) );
  BUFx3_ASAP7_75t_R register___U8655 ( .A(register__n5306), .Y(register__n5305) );
  BUFx2_ASAP7_75t_R register___U8656 ( .A(register__n10798), .Y(register__n5306) );
  BUFx2_ASAP7_75t_R register___U8657 ( .A(register__n5308), .Y(register__n5307) );
  BUFx3_ASAP7_75t_R register___U8658 ( .A(register__n5311), .Y(register__n5310) );
  BUFx2_ASAP7_75t_R register___U8659 ( .A(register__n11164), .Y(register__n5311) );
  BUFx3_ASAP7_75t_R register___U8660 ( .A(register__n11565), .Y(register__n5316) );
  BUFx3_ASAP7_75t_R register___U8661 ( .A(register__n11564), .Y(register__n5317) );
  BUFx3_ASAP7_75t_R register___U8662 ( .A(register__n5320), .Y(register__n5319) );
  BUFx2_ASAP7_75t_R register___U8663 ( .A(register__n11478), .Y(register__n5320) );
  BUFx3_ASAP7_75t_R register___U8664 ( .A(register__n5322), .Y(register__n5321) );
  BUFx2_ASAP7_75t_R register___U8665 ( .A(register__n11477), .Y(register__n5322) );
  INVx2_ASAP7_75t_R register___U8666 ( .A(register__n11476), .Y(register__n5323) );
  BUFx3_ASAP7_75t_R register___U8667 ( .A(register__n5325), .Y(register__n5324) );
  BUFx2_ASAP7_75t_R register___U8668 ( .A(register__n11325), .Y(register__n5325) );
  BUFx3_ASAP7_75t_R register___U8669 ( .A(register__n5327), .Y(register__n5326) );
  BUFx2_ASAP7_75t_R register___U8670 ( .A(register__n7665), .Y(register__n5328) );
  BUFx3_ASAP7_75t_R register___U8671 ( .A(register__n5330), .Y(register__n5329) );
  BUFx2_ASAP7_75t_R register___U8672 ( .A(register__n11324), .Y(register__n5330) );
  BUFx2_ASAP7_75t_R register___U8673 ( .A(register__n9220), .Y(register__n5333) );
  BUFx3_ASAP7_75t_R register___U8674 ( .A(register__n5335), .Y(register__n5334) );
  BUFx2_ASAP7_75t_R register___U8675 ( .A(register__n11199), .Y(register__n5335) );
  BUFx2_ASAP7_75t_R register___U8676 ( .A(register__n11701), .Y(register__n5337) );
  BUFx3_ASAP7_75t_R register___U8677 ( .A(register__n11704), .Y(register__n5338) );
  BUFx3_ASAP7_75t_R register___U8678 ( .A(register__n11703), .Y(register__n5339) );
  BUFx2_ASAP7_75t_R register___U8679 ( .A(register__n8322), .Y(register__n5340) );
  BUFx6f_ASAP7_75t_R register___U8680 ( .A(register__n8247), .Y(register__n12181) );
  BUFx12f_ASAP7_75t_R register___U8681 ( .A(register__n4748), .Y(register__n12182) );
  BUFx12f_ASAP7_75t_R register___U8682 ( .A(register__n5042), .Y(register__n12180) );
  BUFx12f_ASAP7_75t_R register___U8683 ( .A(register__net123601), .Y(register__net64782) );
  BUFx12f_ASAP7_75t_R register___U8684 ( .A(register__n5343), .Y(register__n5342) );
  BUFx12f_ASAP7_75t_R register___U8685 ( .A(register__n3415), .Y(register__n11866) );
  BUFx12f_ASAP7_75t_R register___U8686 ( .A(register__n3544), .Y(register__n5345) );
  BUFx12f_ASAP7_75t_R register___U8687 ( .A(register__n3383), .Y(register__n5346) );
  BUFx12f_ASAP7_75t_R register___U8688 ( .A(register__n3423), .Y(register__n5347) );
  BUFx3_ASAP7_75t_R register___U8689 ( .A(register__net117918), .Y(register__net122533) );
  BUFx12f_ASAP7_75t_R register___U8690 ( .A(register__n5226), .Y(register__n5352) );
  BUFx12f_ASAP7_75t_R register___U8691 ( .A(register__n7907), .Y(register__n5353) );
  BUFx12f_ASAP7_75t_R register___U8692 ( .A(register__n5225), .Y(register__n12475) );
  INVx3_ASAP7_75t_R register___U8693 ( .A(register__n11943), .Y(register__n11934) );
  BUFx12f_ASAP7_75t_R register___U8694 ( .A(register__net122409), .Y(register__net122408) );
  BUFx12f_ASAP7_75t_R register___U8695 ( .A(register__net63300), .Y(register__net122409) );
  BUFx12f_ASAP7_75t_R register___U8696 ( .A(register__net140284), .Y(register__net63286) );
  BUFx12f_ASAP7_75t_R register___U8697 ( .A(register__net122408), .Y(register__net63274) );
  BUFx12f_ASAP7_75t_R register___U8698 ( .A(register__n3168), .Y(register__n5355) );
  BUFx3_ASAP7_75t_R register___U8699 ( .A(register__n5358), .Y(register__n5357) );
  BUFx2_ASAP7_75t_R register___U8700 ( .A(Reg_data[964]), .Y(register__n5358) );
  BUFx3_ASAP7_75t_R register___U8701 ( .A(register__n5360), .Y(register__n5359) );
  BUFx2_ASAP7_75t_R register___U8702 ( .A(Reg_data[963]), .Y(register__n5360) );
  BUFx3_ASAP7_75t_R register___U8703 ( .A(register__net122350), .Y(register__net122349) );
  BUFx2_ASAP7_75t_R register___U8704 ( .A(Reg_data[921]), .Y(register__net122350) );
  BUFx3_ASAP7_75t_R register___U8705 ( .A(register__n5362), .Y(register__n5361) );
  BUFx2_ASAP7_75t_R register___U8706 ( .A(Reg_data[918]), .Y(register__n5362) );
  BUFx3_ASAP7_75t_R register___U8707 ( .A(register__n5364), .Y(register__n5363) );
  BUFx2_ASAP7_75t_R register___U8708 ( .A(Reg_data[917]), .Y(register__n5364) );
  BUFx3_ASAP7_75t_R register___U8709 ( .A(register__n5366), .Y(register__n5365) );
  BUFx2_ASAP7_75t_R register___U8710 ( .A(Reg_data[456]), .Y(register__n5366) );
  BUFx3_ASAP7_75t_R register___U8711 ( .A(register__net122334), .Y(register__net122333) );
  BUFx2_ASAP7_75t_R register___U8712 ( .A(Reg_data[911]), .Y(register__net122334) );
  BUFx3_ASAP7_75t_R register___U8713 ( .A(register__n5368), .Y(register__n5367) );
  BUFx2_ASAP7_75t_R register___U8714 ( .A(Reg_data[910]), .Y(register__n5368) );
  OA22x2_ASAP7_75t_R register___U8715 ( .A1(register__n12427), .A2(register__n1412), .B1(register__n9810), .B2(register__n1418), 
        .Y(register__n12982) );
  INVx1_ASAP7_75t_R register___U8716 ( .A(register__n4146), .Y(register__n5369) );
  OA22x2_ASAP7_75t_R register___U8717 ( .A1(register__net64664), .A2(register__n1549), .B1(register__n7513), .B2(register__n1518), 
        .Y(register__n12599) );
  OA22x2_ASAP7_75t_R register___U8718 ( .A1(register__n12286), .A2(register__n1416), .B1(register__n7821), .B2(register__n1418), 
        .Y(register__n12991) );
  OA22x2_ASAP7_75t_R register___U8719 ( .A1(register__n12293), .A2(register__n11829), .B1(register__n6945), .B2(register__n1529), 
        .Y(register__n12589) );
  OA22x2_ASAP7_75t_R register___U8720 ( .A1(register__net62676), .A2(register__n3120), .B1(register__n7551), .B2(register__n1544), 
        .Y(register__n12579) );
  OA22x2_ASAP7_75t_R register___U8721 ( .A1(register__n12093), .A2(register__n119), .B1(register__n6961), .B2(register__n1522), 
        .Y(register__n12597) );
  OA22x2_ASAP7_75t_R register___U8722 ( .A1(register__n12227), .A2(register__n892), .B1(register__n8540), .B2(register__n898), 
        .Y(register__n13049) );
  INVx1_ASAP7_75t_R register___U8723 ( .A(register__n3859), .Y(register__n5373) );
  OA22x2_ASAP7_75t_R register___U8724 ( .A1(register__n12434), .A2(register__n119), .B1(register__n8207), .B2(register__n1521), 
        .Y(register__n12582) );
  OA22x2_ASAP7_75t_R register___U8725 ( .A1(register__net63014), .A2(register__n4033), .B1(register__n6606), .B2(register__n11917), .Y(register__n12526) );
  INVx4_ASAP7_75t_R register___U8726 ( .A(register__n12033), .Y(register__n12032) );
  BUFx2_ASAP7_75t_R register___U8727 ( .A(register__n3533), .Y(register__n12266) );
  BUFx12f_ASAP7_75t_R register___U8728 ( .A(register__n3068), .Y(register__n12267) );
  INVx1_ASAP7_75t_R register___U8729 ( .A(register__n3014), .Y(register__n5376) );
  INVx1_ASAP7_75t_R register___U8730 ( .A(register__n3016), .Y(register__n5377) );
  INVx1_ASAP7_75t_R register___U8731 ( .A(register__n3018), .Y(register__n5378) );
  OA22x2_ASAP7_75t_R register___U8732 ( .A1(register__n12205), .A2(register__n113), .B1(register__n9599), .B2(register__n1530), 
        .Y(register__n12592) );
  OA22x2_ASAP7_75t_R register___U8733 ( .A1(register__net63996), .A2(register__n2851), .B1(register__net89409), .B2(
        n2840), .Y(register__n13274) );
  OA22x2_ASAP7_75t_R register___U8734 ( .A1(register__net64944), .A2(register__n107), .B1(register__n8345), .B2(register__n1545), 
        .Y(register__n12602) );
  OA22x2_ASAP7_75t_R register___U8735 ( .A1(register__net64856), .A2(register__n3022), .B1(register__net99940), .B2(
        n1601), .Y(register__n12712) );
  INVx1_ASAP7_75t_R register___U8736 ( .A(register__n12712), .Y(register__n5379) );
  OA22x2_ASAP7_75t_R register___U8737 ( .A1(register__net64934), .A2(register__n2825), .B1(register__n8712), .B2(register__n1572), 
        .Y(register__n12883) );
  OA22x2_ASAP7_75t_R register___U8738 ( .A1(register__n12318), .A2(register__n461), .B1(register__n9991), .B2(register__n469), 
        .Y(register__n12929) );
  OA22x2_ASAP7_75t_R register___U8739 ( .A1(register__n11956), .A2(register__n1416), .B1(register__n8763), .B2(register__n1417), 
        .Y(register__n13008) );
  OA22x2_ASAP7_75t_R register___U8740 ( .A1(register__net64922), .A2(register__n576), .B1(register__n10058), .B2(register__n583), 
        .Y(register__n13234) );
  OA22x2_ASAP7_75t_R register___U8741 ( .A1(register__n11990), .A2(register__n3343), .B1(register__n9292), .B2(register__n11781), 
        .Y(register__n12977) );
  INVx1_ASAP7_75t_R register___U8742 ( .A(register__n2921), .Y(register__n5381) );
  OA22x2_ASAP7_75t_R register___U8743 ( .A1(register__net64684), .A2(register__n1974), .B1(register__n10183), .B2(register__n2846), .Y(register__n12911) );
  OA22x2_ASAP7_75t_R register___U8744 ( .A1(register__n12120), .A2(register__n1069), .B1(register__n10229), .B2(register__n81), 
        .Y(register__n12819) );
  OA22x2_ASAP7_75t_R register___U8745 ( .A1(register__n12290), .A2(register__n339), .B1(register__n9820), .B2(register__n68), .Y(
        n12728) );
  OA22x2_ASAP7_75t_R register___U8746 ( .A1(register__net64414), .A2(register__n699), .B1(register__net88817), .B2(register__n685), .Y(register__n13325) );
  OA22x2_ASAP7_75t_R register___U8747 ( .A1(register__n12080), .A2(register__n11730), .B1(register__n10401), .B2(register__n1164), 
        .Y(register__n13380) );
  INVx1_ASAP7_75t_R register___U8748 ( .A(register__n3464), .Y(register__n5386) );
  OA22x2_ASAP7_75t_R register___U8749 ( .A1(register__net62992), .A2(register__n1755), .B1(register__n8813), .B2(register__n3821), 
        .Y(register__n13120) );
  INVx1_ASAP7_75t_R register___U8750 ( .A(register__n3293), .Y(register__n5387) );
  OA22x2_ASAP7_75t_R register___U8751 ( .A1(register__net63006), .A2(register__n1416), .B1(register__n8815), .B2(register__n1419), 
        .Y(register__n12983) );
  OA22x2_ASAP7_75t_R register___U8752 ( .A1(register__n12254), .A2(register__n953), .B1(register__n9646), .B2(register__n958), 
        .Y(register__n13021) );
  INVx2_ASAP7_75t_R register___U8753 ( .A(register__n9485), .Y(register__n10531) );
  INVx2_ASAP7_75t_R register___U8754 ( .A(register__n9547), .Y(register__n11021) );
  INVx2_ASAP7_75t_R register___U8755 ( .A(register__n9491), .Y(register__n10915) );
  INVx2_ASAP7_75t_R register___U8756 ( .A(register__n10347), .Y(register__n10663) );
  BUFx2_ASAP7_75t_R register___U8757 ( .A(register__n11586), .Y(register__n5389) );
  INVx2_ASAP7_75t_R register___U8758 ( .A(register__n9533), .Y(register__n11584) );
  BUFx3_ASAP7_75t_R register___U8759 ( .A(register__n5391), .Y(register__n5390) );
  BUFx2_ASAP7_75t_R register___U8760 ( .A(register__n11442), .Y(register__n5391) );
  BUFx3_ASAP7_75t_R register___U8761 ( .A(register__n5393), .Y(register__n5392) );
  BUFx2_ASAP7_75t_R register___U8762 ( .A(register__n11335), .Y(register__n5393) );
  BUFx2_ASAP7_75t_R register___U8763 ( .A(register__n9171), .Y(register__n5394) );
  BUFx3_ASAP7_75t_R register___U8764 ( .A(register__n5396), .Y(register__n5395) );
  BUFx2_ASAP7_75t_R register___U8765 ( .A(register__n11213), .Y(register__n5396) );
  BUFx3_ASAP7_75t_R register___U8766 ( .A(register__n5398), .Y(register__n5397) );
  BUFx2_ASAP7_75t_R register___U8767 ( .A(register__n10585), .Y(register__n5398) );
  BUFx3_ASAP7_75t_R register___U8768 ( .A(register__n5400), .Y(register__n5399) );
  BUFx2_ASAP7_75t_R register___U8769 ( .A(register__n11466), .Y(register__n5400) );
  BUFx3_ASAP7_75t_R register___U8770 ( .A(register__n5402), .Y(register__n5401) );
  BUFx2_ASAP7_75t_R register___U8771 ( .A(register__n11672), .Y(register__n5402) );
  BUFx2_ASAP7_75t_R register___U8772 ( .A(register__n5404), .Y(register__n5403) );
  BUFx2_ASAP7_75t_R register___U8773 ( .A(register__n12535), .Y(register__n5404) );
  BUFx2_ASAP7_75t_R register___U8774 ( .A(register__n5406), .Y(register__n5405) );
  BUFx2_ASAP7_75t_R register___U8775 ( .A(register__n11188), .Y(register__n5410) );
  BUFx3_ASAP7_75t_R register___U8776 ( .A(register__n5412), .Y(register__n5411) );
  BUFx2_ASAP7_75t_R register___U8777 ( .A(register__n11191), .Y(register__n5412) );
  BUFx3_ASAP7_75t_R register___U8778 ( .A(register__n5417), .Y(register__n5416) );
  BUFx2_ASAP7_75t_R register___U8779 ( .A(register__n10711), .Y(register__n5417) );
  BUFx3_ASAP7_75t_R register___U8780 ( .A(register__n5419), .Y(register__n5418) );
  BUFx2_ASAP7_75t_R register___U8781 ( .A(register__n10709), .Y(register__n5419) );
  BUFx3_ASAP7_75t_R register___U8782 ( .A(register__n5421), .Y(register__n5420) );
  BUFx2_ASAP7_75t_R register___U8783 ( .A(register__n10708), .Y(register__n5421) );
  BUFx2_ASAP7_75t_R register___U8784 ( .A(register__n9151), .Y(register__n5422) );
  BUFx3_ASAP7_75t_R register___U8785 ( .A(register__n5424), .Y(register__n5423) );
  BUFx3_ASAP7_75t_R register___U8786 ( .A(register__n5428), .Y(register__n5427) );
  BUFx2_ASAP7_75t_R register___U8787 ( .A(register__n11423), .Y(register__n5428) );
  BUFx2_ASAP7_75t_R register___U8788 ( .A(register__n6157), .Y(register__n5429) );
  BUFx3_ASAP7_75t_R register___U8789 ( .A(register__n5431), .Y(register__n5430) );
  BUFx2_ASAP7_75t_R register___U8790 ( .A(register__n11378), .Y(register__n5431) );
  BUFx3_ASAP7_75t_R register___U8791 ( .A(register__n5433), .Y(register__n5432) );
  BUFx2_ASAP7_75t_R register___U8792 ( .A(register__n11379), .Y(register__n5433) );
  BUFx3_ASAP7_75t_R register___U8793 ( .A(register__n5438), .Y(register__n5437) );
  BUFx2_ASAP7_75t_R register___U8794 ( .A(register__n11315), .Y(register__n5438) );
  BUFx3_ASAP7_75t_R register___U8795 ( .A(register__n5440), .Y(register__n5439) );
  BUFx2_ASAP7_75t_R register___U8796 ( .A(register__n11312), .Y(register__n5440) );
  BUFx4f_ASAP7_75t_R register___U8797 ( .A(register__n3188), .Y(register__n9405) );
  BUFx6f_ASAP7_75t_R register___U8798 ( .A(register__n3724), .Y(register__n12221) );
  BUFx12f_ASAP7_75t_R register___U8799 ( .A(register__net140664), .Y(register__net121483) );
  BUFx4f_ASAP7_75t_R register___U8800 ( .A(register__net141519), .Y(register__net121484) );
  BUFx12f_ASAP7_75t_R register___U8801 ( .A(register__net100796), .Y(register__net121464) );
  BUFx12f_ASAP7_75t_R register___U8802 ( .A(register__net142807), .Y(register__net62696) );
  BUFx3_ASAP7_75t_R register___U8803 ( .A(register__n5445), .Y(register__n5444) );
  BUFx2_ASAP7_75t_R register___U8804 ( .A(register__n11284), .Y(register__n5445) );
  BUFx2_ASAP7_75t_R register___U8805 ( .A(register__n9234), .Y(register__n5446) );
  BUFx3_ASAP7_75t_R register___U8806 ( .A(register__n5448), .Y(register__n5447) );
  BUFx2_ASAP7_75t_R register___U8807 ( .A(register__n11283), .Y(register__n5448) );
  BUFx3_ASAP7_75t_R register___U8808 ( .A(register__n5450), .Y(register__n5449) );
  BUFx2_ASAP7_75t_R register___U8809 ( .A(register__n11224), .Y(register__n5450) );
  BUFx4f_ASAP7_75t_R register___U8810 ( .A(register__n11222), .Y(register__n8691) );
  INVx2_ASAP7_75t_R register___U8811 ( .A(register__n8691), .Y(register__n5451) );
  BUFx3_ASAP7_75t_R register___U8812 ( .A(register__n5453), .Y(register__n5452) );
  BUFx2_ASAP7_75t_R register___U8813 ( .A(register__n11223), .Y(register__n5453) );
  BUFx2_ASAP7_75t_R register___U8814 ( .A(register__n10951), .Y(register__n5454) );
  BUFx3_ASAP7_75t_R register___U8815 ( .A(register__n5456), .Y(register__n5455) );
  BUFx2_ASAP7_75t_R register___U8816 ( .A(register__n10954), .Y(register__n5456) );
  BUFx2_ASAP7_75t_R register___U8817 ( .A(register__n10953), .Y(register__n5457) );
  BUFx2_ASAP7_75t_R register___U8818 ( .A(register__n10552), .Y(register__n5459) );
  BUFx2_ASAP7_75t_R register___U8819 ( .A(register__n10681), .Y(register__n5460) );
  BUFx3_ASAP7_75t_R register___U8820 ( .A(register__n5463), .Y(register__n5462) );
  BUFx2_ASAP7_75t_R register___U8821 ( .A(register__n10889), .Y(register__n5463) );
  BUFx3_ASAP7_75t_R register___U8822 ( .A(register__n5465), .Y(register__n5464) );
  BUFx2_ASAP7_75t_R register___U8823 ( .A(register__n10888), .Y(register__n5465) );
  BUFx2_ASAP7_75t_R register___U8824 ( .A(register__n8294), .Y(register__n5466) );
  BUFx3_ASAP7_75t_R register___U8825 ( .A(register__n5468), .Y(register__n5467) );
  BUFx2_ASAP7_75t_R register___U8826 ( .A(register__n10738), .Y(register__n5468) );
  BUFx2_ASAP7_75t_R register___U8827 ( .A(register__n10736), .Y(register__n5469) );
  BUFx2_ASAP7_75t_R register___U8828 ( .A(register__n8319), .Y(register__n5470) );
  BUFx3_ASAP7_75t_R register___U8829 ( .A(register__n5475), .Y(register__n5474) );
  BUFx3_ASAP7_75t_R register___U8830 ( .A(register__n5477), .Y(register__n5476) );
  BUFx3_ASAP7_75t_R register___U8831 ( .A(register__n5479), .Y(register__n5478) );
  BUFx2_ASAP7_75t_R register___U8832 ( .A(register__n11683), .Y(register__n5479) );
  BUFx3_ASAP7_75t_R register___U8833 ( .A(register__n5481), .Y(register__n5480) );
  BUFx2_ASAP7_75t_R register___U8834 ( .A(register__n11682), .Y(register__n5481) );
  BUFx3_ASAP7_75t_R register___U8835 ( .A(register__n5483), .Y(register__n5482) );
  BUFx2_ASAP7_75t_R register___U8836 ( .A(register__n11040), .Y(register__n5483) );
  BUFx3_ASAP7_75t_R register___U8837 ( .A(register__n5485), .Y(register__n5484) );
  BUFx2_ASAP7_75t_R register___U8838 ( .A(register__n11039), .Y(register__n5485) );
  BUFx3_ASAP7_75t_R register___U8839 ( .A(register__n5487), .Y(register__n5486) );
  BUFx2_ASAP7_75t_R register___U8840 ( .A(register__n11038), .Y(register__n5487) );
  BUFx2_ASAP7_75t_R register___U8841 ( .A(register__n9205), .Y(register__n5488) );
  BUFx3_ASAP7_75t_R register___U8842 ( .A(register__n5490), .Y(register__n5489) );
  BUFx2_ASAP7_75t_R register___U8843 ( .A(register__n11084), .Y(register__n5490) );
  BUFx3_ASAP7_75t_R register___U8844 ( .A(register__n5492), .Y(register__n5491) );
  BUFx2_ASAP7_75t_R register___U8845 ( .A(register__n11083), .Y(register__n5492) );
  BUFx2_ASAP7_75t_R register___U8846 ( .A(register__n8298), .Y(register__n5493) );
  OR2x2_ASAP7_75t_R register___U8847 ( .A(register__n5496), .B(register__n5495), .Y(register__n5494) );
  BUFx2_ASAP7_75t_R register___U8848 ( .A(register__n8601), .Y(register__n5495) );
  BUFx2_ASAP7_75t_R register___U8849 ( .A(register__n8600), .Y(register__n5496) );
  BUFx12f_ASAP7_75t_R register___U8850 ( .A(register__n12334), .Y(register__n5497) );
  BUFx12f_ASAP7_75t_R register___U8851 ( .A(register__n5347), .Y(register__n12354) );
  BUFx12f_ASAP7_75t_R register___U8852 ( .A(register__n5346), .Y(register__n12351) );
  BUFx12f_ASAP7_75t_R register___U8853 ( .A(register__n5499), .Y(register__n5498) );
  BUFx12f_ASAP7_75t_R register___U8854 ( .A(register__n5504), .Y(register__n5502) );
  BUFx12f_ASAP7_75t_R register___U8855 ( .A(register__n3452), .Y(register__n5503) );
  BUFx12f_ASAP7_75t_R register___U8856 ( .A(register__n3149), .Y(register__n12160) );
  BUFx12f_ASAP7_75t_R register___U8857 ( .A(register__n3044), .Y(register__n12156) );
  BUFx3_ASAP7_75t_R register___U8858 ( .A(register__n7152), .Y(register__n5505) );
  BUFx6f_ASAP7_75t_R register___U8859 ( .A(register__n7151), .Y(register__n9627) );
  BUFx4f_ASAP7_75t_R register___U8860 ( .A(register__n5505), .Y(register__n7151) );
  BUFx3_ASAP7_75t_R register___U8861 ( .A(register__n6288), .Y(register__n5506) );
  BUFx3_ASAP7_75t_R register___U8862 ( .A(register__n5661), .Y(register__n5507) );
  BUFx3_ASAP7_75t_R register___U8863 ( .A(register__n5839), .Y(register__n5508) );
  BUFx3_ASAP7_75t_R register___U8864 ( .A(register__n5840), .Y(register__n5509) );
  BUFx3_ASAP7_75t_R register___U8865 ( .A(register__n6052), .Y(register__n5510) );
  BUFx3_ASAP7_75t_R register___U8866 ( .A(register__n7387), .Y(register__n5511) );
  BUFx3_ASAP7_75t_R register___U8867 ( .A(register__n6054), .Y(register__n5512) );
  BUFx3_ASAP7_75t_R register___U8868 ( .A(register__n7570), .Y(register__n5513) );
  BUFx6f_ASAP7_75t_R register___U8869 ( .A(register__n7569), .Y(register__n8353) );
  BUFx4f_ASAP7_75t_R register___U8870 ( .A(register__n5513), .Y(register__n7569) );
  INVx1_ASAP7_75t_R register___U8871 ( .A(register__n4491), .Y(register__n5517) );
  INVx1_ASAP7_75t_R register___U8872 ( .A(register__n5059), .Y(register__n5518) );
  BUFx12f_ASAP7_75t_R register___U8873 ( .A(register__n3505), .Y(register__n5524) );
  BUFx12f_ASAP7_75t_R register___U8874 ( .A(register__n3506), .Y(register__n5525) );
  BUFx12f_ASAP7_75t_R register___U8875 ( .A(register__n11913), .Y(register__n11836) );
  BUFx3_ASAP7_75t_R register___U8876 ( .A(register__n5527), .Y(register__n5526) );
  BUFx2_ASAP7_75t_R register___U8877 ( .A(Reg_data[644]), .Y(register__n5527) );
  BUFx3_ASAP7_75t_R register___U8878 ( .A(register__n5529), .Y(register__n5528) );
  BUFx2_ASAP7_75t_R register___U8879 ( .A(Reg_data[990]), .Y(register__n5529) );
  INVx2_ASAP7_75t_R register___U8880 ( .A(register__net64790), .Y(register__net64758) );
  BUFx12f_ASAP7_75t_R register___U8881 ( .A(register__n3351), .Y(register__n5530) );
  BUFx12f_ASAP7_75t_R register___U8882 ( .A(register__n3476), .Y(register__n11759) );
  INVx2_ASAP7_75t_R register___U8883 ( .A(register__net91923), .Y(register__net64946) );
  INVx1_ASAP7_75t_R register___U8884 ( .A(register__n11008), .Y(register__n5533) );
  INVx1_ASAP7_75t_R register___U8885 ( .A(register__n3864), .Y(register__n5534) );
  INVx1_ASAP7_75t_R register___U8886 ( .A(register__n4257), .Y(register__n5535) );
  INVx1_ASAP7_75t_R register___U8887 ( .A(register__n4259), .Y(register__n5536) );
  INVx1_ASAP7_75t_R register___U8888 ( .A(register__n4261), .Y(register__n5537) );
  INVx1_ASAP7_75t_R register___U8889 ( .A(register__n2901), .Y(register__n5538) );
  BUFx6f_ASAP7_75t_R register___U8890 ( .A(register__net129902), .Y(register__net64048) );
  BUFx6f_ASAP7_75t_R register___U8891 ( .A(register__net64044), .Y(register__net64042) );
  OA22x2_ASAP7_75t_R register___U8892 ( .A1(register__net63004), .A2(register__n1069), .B1(register__n7220), .B2(register__n3076), 
        .Y(register__n12804) );
  INVx1_ASAP7_75t_R register___U8893 ( .A(register__n3199), .Y(register__n5539) );
  OA22x2_ASAP7_75t_R register___U8894 ( .A1(register__n12032), .A2(register__n4033), .B1(register__n8755), .B2(register__n3216), 
        .Y(register__n12549) );
  OA22x2_ASAP7_75t_R register___U8895 ( .A1(register__n12341), .A2(register__n1569), .B1(register__n8716), .B2(register__n1191), 
        .Y(register__n13094) );
  OA22x2_ASAP7_75t_R register___U8896 ( .A1(register__n12232), .A2(register__n2802), .B1(register__n6778), .B2(register__n1935), 
        .Y(register__n12872) );
  INVx1_ASAP7_75t_R register___U8897 ( .A(register__n3583), .Y(register__n5541) );
  OA22x2_ASAP7_75t_R register___U8898 ( .A1(register__net64670), .A2(register__n578), .B1(register__n10162), .B2(register__n589), 
        .Y(register__n13231) );
  INVx1_ASAP7_75t_R register___U8899 ( .A(register__n3826), .Y(register__n5542) );
  OA22x2_ASAP7_75t_R register___U8900 ( .A1(register__n12091), .A2(register__n3022), .B1(register__n7330), .B2(register__n1605), 
        .Y(register__n12709) );
  OA22x2_ASAP7_75t_R register___U8901 ( .A1(register__net63250), .A2(register__n3343), .B1(register__net93717), .B2(
        n11778), .Y(register__n12955) );
  OA22x2_ASAP7_75t_R register___U8902 ( .A1(register__n12287), .A2(register__n462), .B1(register__n10245), .B2(register__n471), 
        .Y(register__n12930) );
  INVx1_ASAP7_75t_R register___U8903 ( .A(register__n3973), .Y(register__n5544) );
  OA22x2_ASAP7_75t_R register___U8904 ( .A1(register__n12081), .A2(register__n700), .B1(register__n10403), .B2(register__n668), 
        .Y(register__n13326) );
  OA22x2_ASAP7_75t_R register___U8905 ( .A1(register__n12090), .A2(register__n339), .B1(register__n9863), .B2(register__n344), 
        .Y(register__n12738) );
  INVx1_ASAP7_75t_R register___U8906 ( .A(register__n3615), .Y(register__n5545) );
  OA22x2_ASAP7_75t_R register___U8907 ( .A1(register__n12394), .A2(register__n3719), .B1(register__n10405), .B2(register__n1162), 
        .Y(register__n13363) );
  OA22x2_ASAP7_75t_R register___U8908 ( .A1(register__n12170), .A2(register__n890), .B1(register__n9905), .B2(register__n896), 
        .Y(register__n13052) );
  OA22x2_ASAP7_75t_R register___U8909 ( .A1(register__n12171), .A2(register__n1413), .B1(register__n9911), .B2(register__n1418), 
        .Y(register__n12996) );
  INVx1_ASAP7_75t_R register___U8910 ( .A(register__n3589), .Y(register__n5546) );
  OA22x2_ASAP7_75t_R register___U8911 ( .A1(register__n12376), .A2(register__n1755), .B1(register__n9682), .B2(register__n3821), 
        .Y(register__n13125) );
  INVx2_ASAP7_75t_R register___U8912 ( .A(register__n8825), .Y(register__n10960) );
  INVx2_ASAP7_75t_R register___U8913 ( .A(register__n9437), .Y(register__n10826) );
  INVx2_ASAP7_75t_R register___U8914 ( .A(register__n10341), .Y(register__n11247) );
  INVx2_ASAP7_75t_R register___U8915 ( .A(register__n9443), .Y(register__n11205) );
  INVx2_ASAP7_75t_R register___U8916 ( .A(register__n9375), .Y(register__n11183) );
  INVx2_ASAP7_75t_R register___U8917 ( .A(register__n8833), .Y(register__n11353) );
  INVx2_ASAP7_75t_R register___U8918 ( .A(register__n7999), .Y(register__n11503) );
  INVx2_ASAP7_75t_R register___U8919 ( .A(register__n9561), .Y(register__n10789) );
  INVx2_ASAP7_75t_R register___U8920 ( .A(register__n9497), .Y(register__n10599) );
  INVx2_ASAP7_75t_R register___U8921 ( .A(register__n10351), .Y(register__n10556) );
  BUFx2_ASAP7_75t_R register___U8922 ( .A(register__n10663), .Y(register__n5549) );
  BUFx2_ASAP7_75t_R register___U8923 ( .A(register__n10915), .Y(register__n5550) );
  INVx2_ASAP7_75t_R register___U8924 ( .A(register__n10407), .Y(register__n11020) );
  INVx2_ASAP7_75t_R register___U8925 ( .A(register__n9445), .Y(register__n10934) );
  INVx2_ASAP7_75t_R register___U8926 ( .A(register__n9447), .Y(register__n10914) );
  BUFx3_ASAP7_75t_R register___U8927 ( .A(register__n5552), .Y(register__n5551) );
  BUFx2_ASAP7_75t_R register___U8928 ( .A(register__n11574), .Y(register__n5552) );
  BUFx3_ASAP7_75t_R register___U8929 ( .A(register__n5554), .Y(register__n5553) );
  BUFx2_ASAP7_75t_R register___U8930 ( .A(register__n11007), .Y(register__n5554) );
  BUFx3_ASAP7_75t_R register___U8931 ( .A(register__n10630), .Y(register__n5555) );
  BUFx3_ASAP7_75t_R register___U8932 ( .A(register__n5559), .Y(register__n5558) );
  BUFx2_ASAP7_75t_R register___U8933 ( .A(register__n10858), .Y(register__n5559) );
  BUFx3_ASAP7_75t_R register___U8934 ( .A(register__n5561), .Y(register__n5560) );
  BUFx2_ASAP7_75t_R register___U8935 ( .A(register__n10814), .Y(register__n5561) );
  BUFx2_ASAP7_75t_R register___U8936 ( .A(register__n10900), .Y(register__n5562) );
  BUFx2_ASAP7_75t_R register___U8937 ( .A(register__n6300), .Y(register__n5563) );
  BUFx2_ASAP7_75t_R register___U8938 ( .A(register__n5565), .Y(register__n5564) );
  BUFx2_ASAP7_75t_R register___U8939 ( .A(register__n12531), .Y(register__n5565) );
  BUFx2_ASAP7_75t_R register___U8940 ( .A(register__n5567), .Y(register__n5566) );
  BUFx2_ASAP7_75t_R register___U8941 ( .A(register__n12867), .Y(register__n5567) );
  BUFx2_ASAP7_75t_R register___U8942 ( .A(register__n5569), .Y(register__n5568) );
  BUFx2_ASAP7_75t_R register___U8943 ( .A(register__n5571), .Y(register__n5570) );
  BUFx2_ASAP7_75t_R register___U8944 ( .A(register__n5575), .Y(register__n5574) );
  BUFx2_ASAP7_75t_R register___U8945 ( .A(register__n12621), .Y(register__n5575) );
  BUFx2_ASAP7_75t_R register___U8946 ( .A(register__n5577), .Y(register__n5576) );
  BUFx2_ASAP7_75t_R register___U8947 ( .A(register__n12876), .Y(register__n5577) );
  BUFx2_ASAP7_75t_R register___U8948 ( .A(register__n5581), .Y(register__n5580) );
  BUFx2_ASAP7_75t_R register___U8949 ( .A(register__n13210), .Y(register__n5581) );
  BUFx6f_ASAP7_75t_R register___U8950 ( .A(register__n6405), .Y(register__n12011) );
  BUFx3_ASAP7_75t_R register___U8951 ( .A(register__n5583), .Y(register__n5582) );
  BUFx2_ASAP7_75t_R register___U8952 ( .A(register__n10539), .Y(register__n5583) );
  BUFx3_ASAP7_75t_R register___U8953 ( .A(register__n10567), .Y(register__n5584) );
  AO22x1_ASAP7_75t_R register___U8954 ( .A1(register__n5197), .A2(register__n1771), .B1(register__n4180), .B2(register__net126625), .Y(register__n10566) );
  BUFx3_ASAP7_75t_R register___U8955 ( .A(register__n10776), .Y(register__n5585) );
  BUFx3_ASAP7_75t_R register___U8956 ( .A(register__n5590), .Y(register__n5589) );
  BUFx2_ASAP7_75t_R register___U8957 ( .A(register__n11395), .Y(register__n5590) );
  BUFx3_ASAP7_75t_R register___U8958 ( .A(register__n5592), .Y(register__n5591) );
  BUFx2_ASAP7_75t_R register___U8959 ( .A(register__n10695), .Y(register__n5592) );
  BUFx3_ASAP7_75t_R register___U8960 ( .A(register__n5594), .Y(register__n5593) );
  BUFx2_ASAP7_75t_R register___U8961 ( .A(register__n10693), .Y(register__n5594) );
  BUFx3_ASAP7_75t_R register___U8962 ( .A(register__n5596), .Y(register__n5595) );
  BUFx2_ASAP7_75t_R register___U8963 ( .A(register__n10694), .Y(register__n5596) );
  BUFx3_ASAP7_75t_R register___U8964 ( .A(register__n5602), .Y(register__n5601) );
  BUFx2_ASAP7_75t_R register___U8965 ( .A(register__n11692), .Y(register__n5602) );
  BUFx2_ASAP7_75t_R register___U8966 ( .A(register__n6710), .Y(register__n5605) );
  AO22x1_ASAP7_75t_R register___U8967 ( .A1(register__n9796), .A2(register__C6423_net61343), .B1(register__n10116), 
        .B2(register__net122313), .Y(register__n11692) );
  AO22x1_ASAP7_75t_R register___U8968 ( .A1(register__n9788), .A2(register__C6423_net61340), .B1(register__n10104), 
        .B2(register__net125365), .Y(register__n11693) );
  BUFx3_ASAP7_75t_R register___U8969 ( .A(register__n5608), .Y(register__n5607) );
  BUFx2_ASAP7_75t_R register___U8970 ( .A(register__n11296), .Y(register__n5608) );
  BUFx3_ASAP7_75t_R register___U8971 ( .A(register__n5610), .Y(register__n5609) );
  BUFx2_ASAP7_75t_R register___U8972 ( .A(register__n11293), .Y(register__n5610) );
  BUFx3_ASAP7_75t_R register___U8973 ( .A(register__n5614), .Y(register__n5613) );
  BUFx2_ASAP7_75t_R register___U8974 ( .A(register__n11173), .Y(register__n5614) );
  BUFx2_ASAP7_75t_R register___U8975 ( .A(register__n11170), .Y(register__n5615) );
  BUFx3_ASAP7_75t_R register___U8976 ( .A(register__n5620), .Y(register__n5619) );
  BUFx2_ASAP7_75t_R register___U8977 ( .A(register__n11417), .Y(register__n5620) );
  BUFx3_ASAP7_75t_R register___U8978 ( .A(register__n5622), .Y(register__n5621) );
  BUFx2_ASAP7_75t_R register___U8979 ( .A(register__n11416), .Y(register__n5622) );
  BUFx3_ASAP7_75t_R register___U8980 ( .A(register__n5624), .Y(register__n5623) );
  BUFx2_ASAP7_75t_R register___U8981 ( .A(register__n11484), .Y(register__n5624) );
  BUFx2_ASAP7_75t_R register___U8982 ( .A(register__n7948), .Y(register__n5627) );
  BUFx3_ASAP7_75t_R register___U8983 ( .A(register__n10836), .Y(register__n5628) );
  BUFx2_ASAP7_75t_R register___U8984 ( .A(register__n9181), .Y(register__n5629) );
  BUFx12f_ASAP7_75t_R register___U8985 ( .A(register__n7906), .Y(register__n12243) );
  BUFx3_ASAP7_75t_R register___U8986 ( .A(register__n5631), .Y(register__n5630) );
  BUFx2_ASAP7_75t_R register___U8987 ( .A(register__n10978), .Y(register__n5631) );
  BUFx3_ASAP7_75t_R register___U8988 ( .A(register__n5633), .Y(register__n5632) );
  BUFx2_ASAP7_75t_R register___U8989 ( .A(register__n11605), .Y(register__n5633) );
  BUFx3_ASAP7_75t_R register___U8990 ( .A(register__n5635), .Y(register__n5634) );
  BUFx2_ASAP7_75t_R register___U8991 ( .A(register__n11604), .Y(register__n5635) );
  INVx2_ASAP7_75t_R register___U8992 ( .A(register__n11603), .Y(register__n5636) );
  OR2x2_ASAP7_75t_R register___U8993 ( .A(register__n5638), .B(register__n5639), .Y(register__n5637) );
  BUFx2_ASAP7_75t_R register___U8994 ( .A(register__n8661), .Y(register__n5638) );
  OR2x2_ASAP7_75t_R register___U8995 ( .A(register__n12172), .B(register__n1938), .Y(register__n8662) );
  INVx1_ASAP7_75t_R register___U8996 ( .A(register__n3913), .Y(register__n5639) );
  NOR2x1p5_ASAP7_75t_R register___U8997 ( .A(register__n9527), .B(register__n2809), .Y(register__n8661) );
  BUFx12f_ASAP7_75t_R register___U8998 ( .A(register__n5642), .Y(register__n5641) );
  BUFx12f_ASAP7_75t_R register___U8999 ( .A(register__n3325), .Y(register__n5642) );
  BUFx2_ASAP7_75t_R register___U9000 ( .A(register__n9593), .Y(register__n5643) );
  BUFx3_ASAP7_75t_R register___U9001 ( .A(register__n9593), .Y(register__n5644) );
  BUFx4f_ASAP7_75t_R register___U9002 ( .A(register__n9593), .Y(register__n5645) );
  BUFx3_ASAP7_75t_R register___U9003 ( .A(register__n6047), .Y(register__n5646) );
  BUFx3_ASAP7_75t_R register___U9004 ( .A(register__n6048), .Y(register__n5647) );
  BUFx3_ASAP7_75t_R register___U9005 ( .A(register__net88548), .Y(register__net119537) );
  BUFx2_ASAP7_75t_R register___U9006 ( .A(register__net88548), .Y(register__net119539) );
  BUFx3_ASAP7_75t_R register___U9007 ( .A(register__n10001), .Y(register__n5648) );
  BUFx4f_ASAP7_75t_R register___U9008 ( .A(register__n10001), .Y(register__n5649) );
  BUFx2_ASAP7_75t_R register___U9009 ( .A(register__n10001), .Y(register__n5650) );
  BUFx3_ASAP7_75t_R register___U9010 ( .A(register__n6049), .Y(register__n5651) );
  BUFx3_ASAP7_75t_R register___U9011 ( .A(register__n7772), .Y(register__n5652) );
  BUFx6f_ASAP7_75t_R register___U9012 ( .A(register__n7771), .Y(register__n10090) );
  BUFx4f_ASAP7_75t_R register___U9013 ( .A(register__n5652), .Y(register__n7771) );
  BUFx6f_ASAP7_75t_R register___U9014 ( .A(register__n6779), .Y(register__n6778) );
  BUFx3_ASAP7_75t_R register___U9015 ( .A(register__net117906), .Y(register__net119522) );
  BUFx3_ASAP7_75t_R register___U9016 ( .A(register__n6293), .Y(register__n5653) );
  BUFx3_ASAP7_75t_R register___U9017 ( .A(register__n6544), .Y(register__n5654) );
  BUFx3_ASAP7_75t_R register___U9018 ( .A(register__n6294), .Y(register__n5655) );
  BUFx3_ASAP7_75t_R register___U9019 ( .A(register__n6295), .Y(register__n5656) );
  BUFx3_ASAP7_75t_R register___U9020 ( .A(register__n5841), .Y(register__n5657) );
  BUFx3_ASAP7_75t_R register___U9021 ( .A(register__n8173), .Y(register__n5658) );
  BUFx6f_ASAP7_75t_R register___U9022 ( .A(register__n8172), .Y(register__n10268) );
  BUFx4f_ASAP7_75t_R register___U9023 ( .A(register__n5658), .Y(register__n8172) );
  BUFx6f_ASAP7_75t_R register___U9024 ( .A(register__n8352), .Y(register__n8351) );
  BUFx12f_ASAP7_75t_R register___U9025 ( .A(register__n8780), .Y(register__n5659) );
  BUFx3_ASAP7_75t_R register___U9026 ( .A(register__net105576), .Y(register__net119501) );
  BUFx4f_ASAP7_75t_R register___U9027 ( .A(register__net119501), .Y(register__net89010) );
  BUFx12f_ASAP7_75t_R register___U9028 ( .A(register__n11887), .Y(register__n5660) );
  CKINVDCx10_ASAP7_75t_R register___U9029 ( .A(register__n12081), .Y(register__n7257) );
  BUFx12f_ASAP7_75t_R register___U9030 ( .A(register__n12108), .Y(register__n12098) );
  BUFx2_ASAP7_75t_R register___U9031 ( .A(Reg_data[621]), .Y(register__n5661) );
  BUFx6f_ASAP7_75t_R register___U9032 ( .A(register__n10095), .Y(register__n10094) );
  BUFx4f_ASAP7_75t_R register___U9033 ( .A(register__n5507), .Y(register__n10095) );
  BUFx12f_ASAP7_75t_R register___U9034 ( .A(register__n3281), .Y(register__n12469) );
  BUFx12f_ASAP7_75t_R register___U9035 ( .A(register__n3474), .Y(register__n12476) );
  BUFx12f_ASAP7_75t_R register___U9036 ( .A(register__n5352), .Y(register__n12472) );
  INVx1_ASAP7_75t_R register___U9037 ( .A(register__n5401), .Y(register__n5662) );
  INVx1_ASAP7_75t_R register___U9038 ( .A(register__n4493), .Y(register__n5663) );
  INVx1_ASAP7_75t_R register___U9039 ( .A(register__n5250), .Y(register__n5664) );
  INVx1_ASAP7_75t_R register___U9040 ( .A(register__n11119), .Y(register__n5666) );
  INVx3_ASAP7_75t_R register___U9041 ( .A(register__net64868), .Y(register__net64834) );
  BUFx12f_ASAP7_75t_R register___U9042 ( .A(register__n3324), .Y(register__n11761) );
  BUFx12f_ASAP7_75t_R register___U9043 ( .A(register__n4431), .Y(register__n11763) );
  BUFx12f_ASAP7_75t_R register___U9044 ( .A(register__n4578), .Y(register__n12276) );
  BUFx12f_ASAP7_75t_R register___U9045 ( .A(register__n12276), .Y(register__n12265) );
  BUFx3_ASAP7_75t_R register___U9046 ( .A(register__n5668), .Y(register__n5667) );
  BUFx2_ASAP7_75t_R register___U9047 ( .A(Reg_data[808]), .Y(register__n5668) );
  BUFx3_ASAP7_75t_R register___U9048 ( .A(register__n5670), .Y(register__n5669) );
  BUFx2_ASAP7_75t_R register___U9049 ( .A(Reg_data[756]), .Y(register__n5670) );
  BUFx3_ASAP7_75t_R register___U9050 ( .A(register__n5672), .Y(register__n5671) );
  BUFx2_ASAP7_75t_R register___U9051 ( .A(Reg_data[515]), .Y(register__n5672) );
  BUFx3_ASAP7_75t_R register___U9052 ( .A(register__n5674), .Y(register__n5673) );
  BUFx2_ASAP7_75t_R register___U9053 ( .A(Reg_data[212]), .Y(register__n5674) );
  BUFx3_ASAP7_75t_R register___U9054 ( .A(register__n5676), .Y(register__n5675) );
  BUFx2_ASAP7_75t_R register___U9055 ( .A(Reg_data[639]), .Y(register__n5676) );
  BUFx3_ASAP7_75t_R register___U9056 ( .A(register__net119331), .Y(register__net119330) );
  BUFx2_ASAP7_75t_R register___U9057 ( .A(Reg_data[989]), .Y(register__net119331) );
  BUFx3_ASAP7_75t_R register___U9058 ( .A(register__net119327), .Y(register__net119326) );
  BUFx2_ASAP7_75t_R register___U9059 ( .A(Reg_data[527]), .Y(register__net119327) );
  BUFx3_ASAP7_75t_R register___U9060 ( .A(register__n5678), .Y(register__n5677) );
  BUFx2_ASAP7_75t_R register___U9061 ( .A(Reg_data[711]), .Y(register__n5678) );
  BUFx2_ASAP7_75t_R register___U9062 ( .A(register__n10189), .Y(register__n5679) );
  BUFx2_ASAP7_75t_R register___U9063 ( .A(register__n10189), .Y(register__n5680) );
  BUFx4f_ASAP7_75t_R register___U9064 ( .A(register__n10189), .Y(register__n5681) );
  BUFx3_ASAP7_75t_R register___U9065 ( .A(register__n5683), .Y(register__n5682) );
  BUFx2_ASAP7_75t_R register___U9066 ( .A(Reg_data[211]), .Y(register__n5683) );
  INVx2_ASAP7_75t_R register___U9067 ( .A(register__n12208), .Y(register__n12193) );
  BUFx4f_ASAP7_75t_R register___U9068 ( .A(register__n3470), .Y(register__n12208) );
  BUFx12f_ASAP7_75t_R register___U9069 ( .A(register__n5442), .Y(register__n12219) );
  OA22x2_ASAP7_75t_R register___U9070 ( .A1(register__net63158), .A2(register__n577), .B1(register__net89793), .B2(register__n587), .Y(register__n13214) );
  INVx1_ASAP7_75t_R register___U9071 ( .A(register__n3893), .Y(register__n5686) );
  OA22x2_ASAP7_75t_R register___U9072 ( .A1(register__n12322), .A2(register__n11900), .B1(register__n9706), .B2(register__n3262), 
        .Y(register__n12616) );
  OA22x2_ASAP7_75t_R register___U9073 ( .A1(register__n11952), .A2(register__n575), .B1(register__n7466), .B2(register__n580), 
        .Y(register__n13237) );
  INVx1_ASAP7_75t_R register___U9074 ( .A(register__n4517), .Y(register__n5687) );
  INVx1_ASAP7_75t_R register___U9075 ( .A(register__n4108), .Y(register__n5688) );
  INVx1_ASAP7_75t_R register___U9076 ( .A(register__n4110), .Y(register__n5689) );
  INVx1_ASAP7_75t_R register___U9077 ( .A(register__n4113), .Y(register__n5690) );
  AND4x1_ASAP7_75t_R register___U9078 ( .A(register__n5690), .B(register__n5688), .C(register__n6826), .D(register__n4112), .Y(
        n10907) );
  INVx1_ASAP7_75t_R register___U9079 ( .A(register__n4158), .Y(register__n5691) );
  INVx1_ASAP7_75t_R register___U9080 ( .A(register__n4160), .Y(register__n5692) );
  INVx1_ASAP7_75t_R register___U9081 ( .A(register__n4162), .Y(register__n5693) );
  AND4x1_ASAP7_75t_R register___U9082 ( .A(register__n6234), .B(register__n5693), .C(register__n5691), .D(register__n4161), .Y(
        n10860) );
  INVx1_ASAP7_75t_R register___U9083 ( .A(register__n3851), .Y(register__n5694) );
  INVx1_ASAP7_75t_R register___U9084 ( .A(register__n3200), .Y(register__n5695) );
  AO22x2_ASAP7_75t_R register___U9085 ( .A1(register__n6898), .A2(register__n919), .B1(register__n9929), .B2(register__n770), .Y(
        n11577) );
  INVx1_ASAP7_75t_R register___U9086 ( .A(register__n3203), .Y(register__n5696) );
  INVx1_ASAP7_75t_R register___U9087 ( .A(register__n4322), .Y(register__n5697) );
  INVx1_ASAP7_75t_R register___U9088 ( .A(register__n4324), .Y(register__n5698) );
  INVx1_ASAP7_75t_R register___U9089 ( .A(register__n4326), .Y(register__n5699) );
  INVx1_ASAP7_75t_R register___U9090 ( .A(register__n3987), .Y(register__n5700) );
  INVx1_ASAP7_75t_R register___U9091 ( .A(register__n3989), .Y(register__n5701) );
  INVx1_ASAP7_75t_R register___U9092 ( .A(register__n4466), .Y(register__n5704) );
  INVx1_ASAP7_75t_R register___U9093 ( .A(register__n4468), .Y(register__n5705) );
  OA22x2_ASAP7_75t_R register___U9094 ( .A1(register__net63326), .A2(register__n578), .B1(register__n8509), .B2(register__n583), 
        .Y(register__n13215) );
  INVx1_ASAP7_75t_R register___U9095 ( .A(register__n3904), .Y(register__n5707) );
  OA22x2_ASAP7_75t_R register___U9096 ( .A1(register__net64946), .A2(register__n4033), .B1(register__n9254), .B2(register__n11838), .Y(register__n12548) );
  INVx1_ASAP7_75t_R register___U9097 ( .A(register__n3882), .Y(register__n5708) );
  OA22x2_ASAP7_75t_R register___U9098 ( .A1(register__n12348), .A2(register__n110), .B1(register__n7982), .B2(register__n1676), 
        .Y(register__n12642) );
  INVx1_ASAP7_75t_R register___U9099 ( .A(register__n3653), .Y(register__n5709) );
  OA22x2_ASAP7_75t_R register___U9100 ( .A1(register__n11929), .A2(register__n1968), .B1(register__n8714), .B2(register__n2817), 
        .Y(register__n12887) );
  INVx1_ASAP7_75t_R register___U9101 ( .A(register__n3922), .Y(register__n5710) );
  INVx4_ASAP7_75t_R register___U9102 ( .A(register__net64796), .Y(register__net64752) );
  OA22x2_ASAP7_75t_R register___U9103 ( .A1(register__n12021), .A2(register__n575), .B1(register__n10060), .B2(register__n586), 
        .Y(register__n13235) );
  INVx1_ASAP7_75t_R register___U9104 ( .A(register__n4138), .Y(register__n5711) );
  OA22x2_ASAP7_75t_R register___U9105 ( .A1(register__net64344), .A2(register__n461), .B1(register__net89617), .B2(register__n469), .Y(register__n12938) );
  OA22x2_ASAP7_75t_R register___U9106 ( .A1(register__net64340), .A2(register__n891), .B1(register__net90665), .B2(register__n900), .Y(register__n13054) );
  OA22x2_ASAP7_75t_R register___U9107 ( .A1(register__net64350), .A2(register__n575), .B1(register__net89585), .B2(register__n583), .Y(register__n13227) );
  OA22x2_ASAP7_75t_R register___U9108 ( .A1(register__net63998), .A2(register__n578), .B1(register__net96819), .B2(register__n581), .Y(register__n13223) );
  INVx1_ASAP7_75t_R register___U9109 ( .A(register__n4140), .Y(register__n5713) );
  OA22x2_ASAP7_75t_R register___U9110 ( .A1(register__net64006), .A2(register__n101), .B1(register__net93713), .B2(
        n11879), .Y(register__n12964) );
  INVx1_ASAP7_75t_R register___U9111 ( .A(register__n2932), .Y(register__n5714) );
  INVx1_ASAP7_75t_R register___U9112 ( .A(register__n3968), .Y(register__n5715) );
  OA22x2_ASAP7_75t_R register___U9113 ( .A1(register__n12124), .A2(register__n113), .B1(register__n9814), .B2(register__n1537), 
        .Y(register__n12595) );
  OA22x2_ASAP7_75t_R register___U9114 ( .A1(register__n12122), .A2(register__n3022), .B1(register__n7332), .B2(register__n1594), 
        .Y(register__n12706) );
  OA22x2_ASAP7_75t_R register___U9115 ( .A1(register__n12287), .A2(register__n1973), .B1(register__n10469), .B2(register__n11785), 
        .Y(register__n12900) );
  INVx1_ASAP7_75t_R register___U9116 ( .A(register__n3224), .Y(register__n5717) );
  OA22x2_ASAP7_75t_R register___U9117 ( .A1(register__n12111), .A2(register__n702), .B1(register__n10409), .B2(register__n684), 
        .Y(register__n13323) );
  OA22x2_ASAP7_75t_R register___U9118 ( .A1(register__net63258), .A2(register__n115), .B1(register__net89037), .B2(
        n1624), .Y(register__n12753) );
  OA22x2_ASAP7_75t_R register___U9119 ( .A1(register__net62984), .A2(register__n3719), .B1(register__n10411), .B2(register__n1162), .Y(register__n13362) );
  INVx1_ASAP7_75t_R register___U9120 ( .A(register__n2860), .Y(register__n5722) );
  OA22x2_ASAP7_75t_R register___U9121 ( .A1(register__n12340), .A2(register__n1266), .B1(register__n9684), .B2(register__n3821), 
        .Y(register__n13126) );
  OA22x2_ASAP7_75t_R register___U9122 ( .A1(register__n12085), .A2(register__n957), .B1(register__n9730), .B2(register__n958), 
        .Y(register__n13029) );
  INVx2_ASAP7_75t_R register___U9123 ( .A(register__n9435), .Y(register__n10959) );
  INVx2_ASAP7_75t_R register___U9124 ( .A(register__n9481), .Y(register__n10598) );
  BUFx2_ASAP7_75t_R register___U9125 ( .A(register__n10826), .Y(register__n5724) );
  INVx2_ASAP7_75t_R register___U9126 ( .A(register__n10345), .Y(register__n11206) );
  BUFx2_ASAP7_75t_R register___U9127 ( .A(register__n10960), .Y(register__n5725) );
  INVx2_ASAP7_75t_R register___U9128 ( .A(register__n9519), .Y(register__n10642) );
  BUFx2_ASAP7_75t_R register___U9129 ( .A(register__n11352), .Y(register__n5726) );
  BUFx2_ASAP7_75t_R register___U9130 ( .A(register__n10743), .Y(register__n5727) );
  INVx2_ASAP7_75t_R register___U9131 ( .A(register__n10349), .Y(register__n10621) );
  BUFx2_ASAP7_75t_R register___U9132 ( .A(register__n10599), .Y(register__n5730) );
  INVx2_ASAP7_75t_R register___U9133 ( .A(register__n9489), .Y(register__n11547) );
  BUFx2_ASAP7_75t_R register___U9134 ( .A(register__C6422_net59963), .Y(register__net118829) );
  BUFx2_ASAP7_75t_R register___U9135 ( .A(register__n11373), .Y(register__n5731) );
  INVx2_ASAP7_75t_R register___U9136 ( .A(register__n9461), .Y(register__n10935) );
  INVx2_ASAP7_75t_R register___U9137 ( .A(register__n9457), .Y(register__n10530) );
  BUFx2_ASAP7_75t_R register___U9138 ( .A(register__n10979), .Y(register__n5732) );
  BUFx2_ASAP7_75t_R register___U9139 ( .A(register__n11584), .Y(register__n5733) );
  BUFx3_ASAP7_75t_R register___U9140 ( .A(register__n11291), .Y(register__n5736) );
  BUFx3_ASAP7_75t_R register___U9141 ( .A(register__n5738), .Y(register__n5737) );
  BUFx2_ASAP7_75t_R register___U9142 ( .A(register__n11272), .Y(register__n5738) );
  BUFx3_ASAP7_75t_R register___U9143 ( .A(register__n5740), .Y(register__n5739) );
  BUFx2_ASAP7_75t_R register___U9144 ( .A(register__n11230), .Y(register__n5740) );
  AO22x1_ASAP7_75t_R register___U9145 ( .A1(register__n6961), .A2(register__n268), .B1(register__n6625), .B2(
        C6423_net61317), .Y(register__n11356) );
  BUFx3_ASAP7_75t_R register___U9146 ( .A(register__n5746), .Y(register__n5745) );
  BUFx2_ASAP7_75t_R register___U9147 ( .A(register__n5748), .Y(register__n5747) );
  BUFx2_ASAP7_75t_R register___U9148 ( .A(register__n5752), .Y(register__n5751) );
  BUFx2_ASAP7_75t_R register___U9149 ( .A(register__n12945), .Y(register__n5752) );
  BUFx2_ASAP7_75t_R register___U9150 ( .A(register__n5754), .Y(register__n5753) );
  BUFx2_ASAP7_75t_R register___U9151 ( .A(register__n5756), .Y(register__n5755) );
  BUFx2_ASAP7_75t_R register___U9152 ( .A(register__n5758), .Y(register__n5757) );
  BUFx2_ASAP7_75t_R register___U9153 ( .A(register__n13063), .Y(register__n5758) );
  BUFx2_ASAP7_75t_R register___U9154 ( .A(register__n5762), .Y(register__n5761) );
  BUFx2_ASAP7_75t_R register___U9155 ( .A(register__n12628), .Y(register__n5762) );
  BUFx2_ASAP7_75t_R register___U9156 ( .A(register__n5768), .Y(register__n5767) );
  NOR2x2_ASAP7_75t_R register___U9157 ( .A(register__n984), .B(register__net64838), .Y(register__n5769) );
  BUFx2_ASAP7_75t_R register___U9158 ( .A(register__n5772), .Y(register__n5771) );
  BUFx2_ASAP7_75t_R register___U9159 ( .A(register__n12522), .Y(register__n5772) );
  BUFx2_ASAP7_75t_R register___U9160 ( .A(register__n5778), .Y(register__n5777) );
  INVx2_ASAP7_75t_R register___U9161 ( .A(register__n12134), .Y(register__n12118) );
  BUFx2_ASAP7_75t_R register___U9162 ( .A(register__n5782), .Y(register__n5781) );
  INVx6_ASAP7_75t_R register___U9163 ( .A(register__n12470), .Y(register__n12455) );
  BUFx2_ASAP7_75t_R register___U9164 ( .A(register__n12692), .Y(register__n5786) );
  BUFx2_ASAP7_75t_R register___U9165 ( .A(register__n13198), .Y(register__n5788) );
  BUFx2_ASAP7_75t_R register___U9166 ( .A(register__n5790), .Y(register__n5789) );
  BUFx2_ASAP7_75t_R register___U9167 ( .A(register__n12695), .Y(register__n5790) );
  BUFx2_ASAP7_75t_R register___U9168 ( .A(register__n5792), .Y(register__n5791) );
  BUFx2_ASAP7_75t_R register___U9169 ( .A(register__n5794), .Y(register__n5793) );
  BUFx2_ASAP7_75t_R register___U9170 ( .A(register__n13111), .Y(register__n5794) );
  BUFx3_ASAP7_75t_R register___U9171 ( .A(register__n5802), .Y(register__n5801) );
  BUFx2_ASAP7_75t_R register___U9172 ( .A(register__n11169), .Y(register__n5802) );
  BUFx3_ASAP7_75t_R register___U9173 ( .A(register__n5807), .Y(register__n5806) );
  BUFx2_ASAP7_75t_R register___U9174 ( .A(register__n11178), .Y(register__n5807) );
  BUFx3_ASAP7_75t_R register___U9175 ( .A(register__n5809), .Y(register__n5808) );
  BUFx4f_ASAP7_75t_R register___U9176 ( .A(register__n5808), .Y(register__n8745) );
  INVx2_ASAP7_75t_R register___U9177 ( .A(register__n8745), .Y(register__n5810) );
  BUFx3_ASAP7_75t_R register___U9178 ( .A(register__n5812), .Y(register__n5811) );
  BUFx2_ASAP7_75t_R register___U9179 ( .A(register__n11177), .Y(register__n5812) );
  BUFx3_ASAP7_75t_R register___U9180 ( .A(register__n5814), .Y(register__n5813) );
  BUFx3_ASAP7_75t_R register___U9181 ( .A(register__n5816), .Y(register__n5815) );
  BUFx2_ASAP7_75t_R register___U9182 ( .A(register__n11389), .Y(register__n5816) );
  BUFx3_ASAP7_75t_R register___U9183 ( .A(register__n5818), .Y(register__n5817) );
  BUFx2_ASAP7_75t_R register___U9184 ( .A(register__n8705), .Y(register__n5819) );
  BUFx3_ASAP7_75t_R register___U9185 ( .A(register__n5821), .Y(register__n5820) );
  BUFx3_ASAP7_75t_R register___U9186 ( .A(register__n5823), .Y(register__n5822) );
  BUFx2_ASAP7_75t_R register___U9187 ( .A(register__n11410), .Y(register__n5823) );
  BUFx3_ASAP7_75t_R register___U9188 ( .A(register__n5825), .Y(register__n5824) );
  BUFx2_ASAP7_75t_R register___U9189 ( .A(register__n7981), .Y(register__n5827) );
  BUFx3_ASAP7_75t_R register___U9190 ( .A(register__n6287), .Y(register__n5828) );
  BUFx3_ASAP7_75t_R register___U9191 ( .A(register__net106228), .Y(register__net118041) );
  BUFx4f_ASAP7_75t_R register___U9192 ( .A(register__net118041), .Y(register__net97214) );
  BUFx3_ASAP7_75t_R register___U9193 ( .A(register__n8963), .Y(register__n5829) );
  BUFx6f_ASAP7_75t_R register___U9194 ( .A(register__n8962), .Y(register__n10093) );
  BUFx4f_ASAP7_75t_R register___U9195 ( .A(register__n5829), .Y(register__n8962) );
  BUFx3_ASAP7_75t_R register___U9196 ( .A(register__n8088), .Y(register__n5830) );
  BUFx6f_ASAP7_75t_R register___U9197 ( .A(register__n8087), .Y(register__n10462) );
  BUFx4f_ASAP7_75t_R register___U9198 ( .A(register__n5830), .Y(register__n8087) );
  BUFx3_ASAP7_75t_R register___U9199 ( .A(register__n8111), .Y(register__n5831) );
  BUFx3_ASAP7_75t_R register___U9200 ( .A(register__n6053), .Y(register__n5832) );
  BUFx3_ASAP7_75t_R register___U9201 ( .A(register__n9028), .Y(register__n5833) );
  BUFx6f_ASAP7_75t_R register___U9202 ( .A(register__n9027), .Y(register__n10164) );
  BUFx4f_ASAP7_75t_R register___U9203 ( .A(register__n5833), .Y(register__n9027) );
  BUFx3_ASAP7_75t_R register___U9204 ( .A(register__net112592), .Y(register__net118023) );
  BUFx3_ASAP7_75t_R register___U9205 ( .A(register__n9042), .Y(register__n5834) );
  BUFx3_ASAP7_75t_R register___U9206 ( .A(register__n9327), .Y(register__n5835) );
  BUFx2_ASAP7_75t_R register___U9207 ( .A(register__n9327), .Y(register__n5836) );
  BUFx3_ASAP7_75t_R register___U9208 ( .A(register__n6055), .Y(register__n5837) );
  BUFx3_ASAP7_75t_R register___U9209 ( .A(register__net100903), .Y(register__net118011) );
  BUFx12f_ASAP7_75t_R register___U9210 ( .A(register__n6301), .Y(register__n11888) );
  AND3x1_ASAP7_75t_R register___U9211 ( .A(register__n1511), .B(register__n12510), .C(register__n12511), .Y(register__n12509) );
  BUFx2_ASAP7_75t_R register___U9212 ( .A(Reg_data[518]), .Y(register__net117918) );
  BUFx4f_ASAP7_75t_R register___U9213 ( .A(register__net122533), .Y(register__net91563) );
  BUFx2_ASAP7_75t_R register___U9214 ( .A(Reg_data[511]), .Y(register__n5839) );
  BUFx6f_ASAP7_75t_R register___U9215 ( .A(register__n10502), .Y(register__n10501) );
  BUFx4f_ASAP7_75t_R register___U9216 ( .A(register__n5508), .Y(register__n10502) );
  BUFx2_ASAP7_75t_R register___U9217 ( .A(Reg_data[631]), .Y(register__n5840) );
  BUFx6f_ASAP7_75t_R register___U9218 ( .A(register__n10123), .Y(register__n10122) );
  BUFx4f_ASAP7_75t_R register___U9219 ( .A(register__n5509), .Y(register__n10123) );
  BUFx2_ASAP7_75t_R register___U9220 ( .A(Reg_data[47]), .Y(register__net117906) );
  BUFx4f_ASAP7_75t_R register___U9221 ( .A(register__net119522), .Y(register__net89553) );
  BUFx2_ASAP7_75t_R register___U9222 ( .A(Reg_data[407]), .Y(register__n5841) );
  BUFx6f_ASAP7_75t_R register___U9223 ( .A(register__n9416), .Y(register__n9415) );
  BUFx4f_ASAP7_75t_R register___U9224 ( .A(register__n5657), .Y(register__n9416) );
  INVx1_ASAP7_75t_R register___U9225 ( .A(register__n5256), .Y(register__n5842) );
  INVx1_ASAP7_75t_R register___U9226 ( .A(register__n5551), .Y(register__n5844) );
  BUFx3_ASAP7_75t_R register___U9227 ( .A(register__n5846), .Y(register__n5845) );
  BUFx2_ASAP7_75t_R register___U9228 ( .A(Reg_data[982]), .Y(register__n5846) );
  BUFx3_ASAP7_75t_R register___U9229 ( .A(register__n5848), .Y(register__n5847) );
  BUFx2_ASAP7_75t_R register___U9230 ( .A(Reg_data[978]), .Y(register__n5848) );
  BUFx3_ASAP7_75t_R register___U9231 ( .A(register__n5850), .Y(register__n5849) );
  BUFx2_ASAP7_75t_R register___U9232 ( .A(Reg_data[968]), .Y(register__n5850) );
  BUFx3_ASAP7_75t_R register___U9233 ( .A(register__n5852), .Y(register__n5851) );
  BUFx2_ASAP7_75t_R register___U9234 ( .A(Reg_data[961]), .Y(register__n5852) );
  BUFx3_ASAP7_75t_R register___U9235 ( .A(register__n5854), .Y(register__n5853) );
  BUFx2_ASAP7_75t_R register___U9236 ( .A(Reg_data[801]), .Y(register__n5854) );
  BUFx3_ASAP7_75t_R register___U9237 ( .A(register__n5856), .Y(register__n5855) );
  BUFx2_ASAP7_75t_R register___U9238 ( .A(Reg_data[757]), .Y(register__n5856) );
  BUFx3_ASAP7_75t_R register___U9239 ( .A(register__n5858), .Y(register__n5857) );
  BUFx2_ASAP7_75t_R register___U9240 ( .A(Reg_data[754]), .Y(register__n5858) );
  BUFx3_ASAP7_75t_R register___U9241 ( .A(register__n5860), .Y(register__n5859) );
  BUFx2_ASAP7_75t_R register___U9242 ( .A(Reg_data[752]), .Y(register__n5860) );
  BUFx3_ASAP7_75t_R register___U9243 ( .A(register__net117776), .Y(register__net117775) );
  BUFx2_ASAP7_75t_R register___U9244 ( .A(Reg_data[742]), .Y(register__net117776) );
  BUFx3_ASAP7_75t_R register___U9245 ( .A(register__n5862), .Y(register__n5861) );
  BUFx2_ASAP7_75t_R register___U9246 ( .A(Reg_data[706]), .Y(register__n5862) );
  BUFx3_ASAP7_75t_R register___U9247 ( .A(register__n5864), .Y(register__n5863) );
  BUFx2_ASAP7_75t_R register___U9248 ( .A(Reg_data[680]), .Y(register__n5864) );
  BUFx3_ASAP7_75t_R register___U9249 ( .A(register__n5866), .Y(register__n5865) );
  BUFx2_ASAP7_75t_R register___U9250 ( .A(Reg_data[616]), .Y(register__n5866) );
  BUFx3_ASAP7_75t_R register___U9251 ( .A(register__n5868), .Y(register__n5867) );
  BUFx2_ASAP7_75t_R register___U9252 ( .A(Reg_data[533]), .Y(register__n5868) );
  BUFx3_ASAP7_75t_R register___U9253 ( .A(register__n5870), .Y(register__n5869) );
  BUFx2_ASAP7_75t_R register___U9254 ( .A(Reg_data[532]), .Y(register__n5870) );
  BUFx3_ASAP7_75t_R register___U9255 ( .A(register__n5872), .Y(register__n5871) );
  BUFx2_ASAP7_75t_R register___U9256 ( .A(Reg_data[8]), .Y(register__n5872) );
  BUFx3_ASAP7_75t_R register___U9257 ( .A(register__net117748), .Y(register__net117747) );
  BUFx2_ASAP7_75t_R register___U9258 ( .A(Reg_data[6]), .Y(register__net117748) );
  BUFx3_ASAP7_75t_R register___U9259 ( .A(register__n5874), .Y(register__n5873) );
  BUFx2_ASAP7_75t_R register___U9260 ( .A(Reg_data[397]), .Y(register__n5874) );
  BUFx3_ASAP7_75t_R register___U9261 ( .A(register__n5876), .Y(register__n5875) );
  BUFx2_ASAP7_75t_R register___U9262 ( .A(Reg_data[169]), .Y(register__n5876) );
  BUFx3_ASAP7_75t_R register___U9263 ( .A(register__n10173), .Y(register__n5877) );
  BUFx2_ASAP7_75t_R register___U9264 ( .A(register__n10173), .Y(register__n5878) );
  BUFx3_ASAP7_75t_R register___U9265 ( .A(register__n5880), .Y(register__n5879) );
  BUFx2_ASAP7_75t_R register___U9266 ( .A(Reg_data[222]), .Y(register__n5880) );
  BUFx3_ASAP7_75t_R register___U9267 ( .A(register__n5882), .Y(register__n5881) );
  BUFx2_ASAP7_75t_R register___U9268 ( .A(Reg_data[206]), .Y(register__n5882) );
  BUFx3_ASAP7_75t_R register___U9269 ( .A(register__n5884), .Y(register__n5883) );
  BUFx2_ASAP7_75t_R register___U9270 ( .A(Reg_data[254]), .Y(register__n5884) );
  BUFx3_ASAP7_75t_R register___U9271 ( .A(register__n5886), .Y(register__n5885) );
  BUFx2_ASAP7_75t_R register___U9272 ( .A(Reg_data[750]), .Y(register__n5886) );
  BUFx3_ASAP7_75t_R register___U9273 ( .A(register__net117708), .Y(register__net117707) );
  BUFx2_ASAP7_75t_R register___U9274 ( .A(Reg_data[938]), .Y(register__net117708) );
  BUFx2_ASAP7_75t_R register___U9275 ( .A(register__net90453), .Y(register__net117709) );
  BUFx3_ASAP7_75t_R register___U9276 ( .A(register__net90453), .Y(register__net117710) );
  BUFx3_ASAP7_75t_R register___U9277 ( .A(register__n5888), .Y(register__n5887) );
  BUFx2_ASAP7_75t_R register___U9278 ( .A(Reg_data[748]), .Y(register__n5888) );
  BUFx3_ASAP7_75t_R register___U9279 ( .A(register__n5890), .Y(register__n5889) );
  BUFx2_ASAP7_75t_R register___U9280 ( .A(Reg_data[755]), .Y(register__n5890) );
  BUFx3_ASAP7_75t_R register___U9281 ( .A(register__n5892), .Y(register__n5891) );
  BUFx2_ASAP7_75t_R register___U9282 ( .A(Reg_data[735]), .Y(register__n5892) );
  BUFx3_ASAP7_75t_R register___U9283 ( .A(register__n5894), .Y(register__n5893) );
  BUFx2_ASAP7_75t_R register___U9284 ( .A(Reg_data[753]), .Y(register__n5894) );
  BUFx3_ASAP7_75t_R register___U9285 ( .A(register__n5896), .Y(register__n5895) );
  BUFx2_ASAP7_75t_R register___U9286 ( .A(Reg_data[913]), .Y(register__n5896) );
  BUFx12f_ASAP7_75t_R register___U9287 ( .A(register__net121463), .Y(register__net62710) );
  OA22x2_ASAP7_75t_R register___U9288 ( .A1(register__net64916), .A2(register__n11730), .B1(register__n10355), .B2(
        n1164), .Y(register__n13384) );
  INVx1_ASAP7_75t_R register___U9289 ( .A(register__n3951), .Y(register__n5897) );
  INVx6_ASAP7_75t_R register___U9290 ( .A(register__n11968), .Y(register__n11952) );
  OA22x2_ASAP7_75t_R register___U9291 ( .A1(register__n12235), .A2(register__n4267), .B1(register__n9724), .B2(register__n3153), 
        .Y(register__n12619) );
  INVx1_ASAP7_75t_R register___U9292 ( .A(register__n4661), .Y(register__n5900) );
  OA22x2_ASAP7_75t_R register___U9293 ( .A1(register__net64686), .A2(register__n339), .B1(register__n9778), .B2(register__n68), 
        .Y(register__n12740) );
  OA22x2_ASAP7_75t_R register___U9294 ( .A1(register__net62816), .A2(register__n11730), .B1(register__net88764), .B2(
        n1164), .Y(register__n13360) );
  INVx1_ASAP7_75t_R register___U9295 ( .A(register__n4011), .Y(register__n5903) );
  INVx6_ASAP7_75t_R register___U9296 ( .A(register__net141520), .Y(register__net62816) );
  OA22x2_ASAP7_75t_R register___U9297 ( .A1(register__n12348), .A2(register__n4267), .B1(register__n9704), .B2(register__n4841), 
        .Y(register__n12615) );
  INVx1_ASAP7_75t_R register___U9298 ( .A(register__n4511), .Y(register__n5904) );
  OA22x2_ASAP7_75t_R register___U9299 ( .A1(register__n12176), .A2(register__n4267), .B1(register__n9802), .B2(register__n11823), 
        .Y(register__n12622) );
  INVx1_ASAP7_75t_R register___U9300 ( .A(register__n12622), .Y(register__n5905) );
  OA22x2_ASAP7_75t_R register___U9301 ( .A1(register__n12147), .A2(register__n1092), .B1(register__n8106), .B2(register__n4431), 
        .Y(register__n13078) );
  OA22x2_ASAP7_75t_R register___U9302 ( .A1(register__net64004), .A2(register__n890), .B1(register__net114113), .B2(
        n897), .Y(register__n13051) );
  OA22x2_ASAP7_75t_R register___U9303 ( .A1(register__n12172), .A2(register__n460), .B1(register__n6385), .B2(register__n467), 
        .Y(register__n12935) );
  OA22x2_ASAP7_75t_R register___U9304 ( .A1(register__n12404), .A2(register__n337), .B1(register__n9096), .B2(register__n342), 
        .Y(register__n12722) );
  INVx1_ASAP7_75t_R register___U9305 ( .A(register__n4535), .Y(register__n5908) );
  OA22x2_ASAP7_75t_R register___U9306 ( .A1(register__n12399), .A2(register__n894), .B1(register__n9112), .B2(register__n904), 
        .Y(register__n13042) );
  OA22x2_ASAP7_75t_R register___U9307 ( .A1(register__n12231), .A2(register__n459), .B1(register__n7563), .B2(register__n466), 
        .Y(register__n12932) );
  INVx1_ASAP7_75t_R register___U9308 ( .A(register__n3976), .Y(register__n5910) );
  OA22x2_ASAP7_75t_R register___U9309 ( .A1(register__net62832), .A2(register__n459), .B1(register__net98193), .B2(register__n466), .Y(register__n12921) );
  OA22x2_ASAP7_75t_R register___U9310 ( .A1(register__n12116), .A2(register__n889), .B1(register__n8529), .B2(register__n900), 
        .Y(register__n13053) );
  OA22x2_ASAP7_75t_R register___U9311 ( .A1(register__net63010), .A2(register__n11900), .B1(register__n7538), .B2(
        n11903), .Y(register__n12609) );
  INVx1_ASAP7_75t_R register___U9312 ( .A(register__n4554), .Y(register__n5914) );
  AND4x1_ASAP7_75t_R register___U9313 ( .A(register__n5914), .B(register__n1256), .C(register__n1460), .D(register__n4553), .Y(
        n10839) );
  INVx1_ASAP7_75t_R register___U9314 ( .A(register__n5430), .Y(register__n5917) );
  INVx1_ASAP7_75t_R register___U9315 ( .A(register__n5432), .Y(register__n5918) );
  INVx1_ASAP7_75t_R register___U9316 ( .A(register__n5434), .Y(register__n5919) );
  AO22x1_ASAP7_75t_R register___U9317 ( .A1(register__n9605), .A2(register__C6423_net61318), .B1(register__n10030), 
        .B2(register__n1448), .Y(register__n11164) );
  INVx1_ASAP7_75t_R register___U9318 ( .A(register__n5310), .Y(register__n5920) );
  INVx1_ASAP7_75t_R register___U9319 ( .A(register__n4432), .Y(register__n5921) );
  INVx1_ASAP7_75t_R register___U9320 ( .A(register__n4434), .Y(register__n5922) );
  INVx1_ASAP7_75t_R register___U9321 ( .A(register__n4437), .Y(register__n5923) );
  INVx1_ASAP7_75t_R register___U9322 ( .A(register__n5437), .Y(register__n5924) );
  INVx1_ASAP7_75t_R register___U9323 ( .A(register__n5439), .Y(register__n5925) );
  INVx1_ASAP7_75t_R register___U9324 ( .A(register__n11113), .Y(register__n5926) );
  AND4x1_ASAP7_75t_R register___U9325 ( .A(register__n5926), .B(register__n5927), .C(register__n292), .D(register__n4026), .Y(
        n11097) );
  OA22x2_ASAP7_75t_R register___U9326 ( .A1(register__n12375), .A2(register__n4035), .B1(register__n7657), .B2(register__n1590), 
        .Y(register__n12698) );
  INVx1_ASAP7_75t_R register___U9327 ( .A(register__n3855), .Y(register__n5930) );
  OA22x2_ASAP7_75t_R register___U9328 ( .A1(register__net62838), .A2(register__n337), .B1(register__net114504), .B2(
        n346), .Y(register__n12719) );
  OA22x2_ASAP7_75t_R register___U9329 ( .A1(register__net120805), .A2(register__n4033), .B1(register__net91105), .B2(
        n11843), .Y(register__n12546) );
  OA22x2_ASAP7_75t_R register___U9330 ( .A1(register__n11998), .A2(register__n4033), .B1(register__n9575), .B2(register__n11916), 
        .Y(register__n12550) );
  OA22x2_ASAP7_75t_R register___U9331 ( .A1(register__n12322), .A2(register__n2116), .B1(register__n7954), .B2(register__n1666), 
        .Y(register__n12643) );
  INVx1_ASAP7_75t_R register___U9332 ( .A(register__n3682), .Y(register__n5932) );
  OA22x2_ASAP7_75t_R register___U9333 ( .A1(register__n12374), .A2(register__n339), .B1(register__n9621), .B2(register__n343), 
        .Y(register__n12725) );
  INVx1_ASAP7_75t_R register___U9334 ( .A(register__n3573), .Y(register__n5933) );
  OA22x2_ASAP7_75t_R register___U9335 ( .A1(register__n12320), .A2(register__n337), .B1(register__n9623), .B2(register__n346), 
        .Y(register__n12727) );
  INVx1_ASAP7_75t_R register___U9336 ( .A(register__n4495), .Y(register__n5934) );
  OA22x2_ASAP7_75t_R register___U9337 ( .A1(register__net64938), .A2(register__n341), .B1(register__n9628), .B2(register__n344), 
        .Y(register__n12742) );
  OA22x2_ASAP7_75t_R register___U9338 ( .A1(register__n12026), .A2(register__n462), .B1(register__n9995), .B2(register__n472), 
        .Y(register__n12946) );
  INVx1_ASAP7_75t_R register___U9339 ( .A(register__n4775), .Y(register__n5935) );
  OA22x2_ASAP7_75t_R register___U9340 ( .A1(register__net63164), .A2(register__n890), .B1(register__net90877), .B2(register__n898), .Y(register__n13043) );
  OA22x2_ASAP7_75t_R register___U9341 ( .A1(register__n12369), .A2(register__n890), .B1(register__n8765), .B2(register__n901), 
        .Y(register__n13045) );
  INVx1_ASAP7_75t_R register___U9342 ( .A(register__n5077), .Y(register__n5936) );
  OA22x2_ASAP7_75t_R register___U9343 ( .A1(register__net64920), .A2(register__n2834), .B1(register__n10026), .B2(register__n3297), .Y(register__n13281) );
  OA22x2_ASAP7_75t_R register___U9344 ( .A1(register__n12343), .A2(register__n11730), .B1(register__n9503), .B2(register__n1164), 
        .Y(register__n13368) );
  OA22x2_ASAP7_75t_R register___U9345 ( .A1(register__n12146), .A2(register__n1137), .B1(register__n9507), .B2(register__n1144), 
        .Y(register__n13164) );
  INVx1_ASAP7_75t_R register___U9346 ( .A(register__n4078), .Y(register__n5939) );
  INVx4_ASAP7_75t_R register___U9347 ( .A(register__net139861), .Y(register__net64682) );
  OA22x2_ASAP7_75t_R register___U9348 ( .A1(register__net63992), .A2(register__n3719), .B1(register__net91259), .B2(
        n1164), .Y(register__n13374) );
  OA22x2_ASAP7_75t_R register___U9349 ( .A1(register__n12110), .A2(register__n3719), .B1(register__n9553), .B2(register__n1162), 
        .Y(register__n13377) );
  OA22x2_ASAP7_75t_R register___U9350 ( .A1(register__n3501), .A2(register__n100), .B1(register__n9244), .B2(register__n11769), 
        .Y(register__n12976) );
  INVx1_ASAP7_75t_R register___U9351 ( .A(register__n2943), .Y(register__n5940) );
  OA22x2_ASAP7_75t_R register___U9352 ( .A1(register__net129768), .A2(register__n462), .B1(register__n10181), .B2(register__n464), 
        .Y(register__n12942) );
  INVx1_ASAP7_75t_R register___U9353 ( .A(register__n4779), .Y(register__n5941) );
  OA22x2_ASAP7_75t_R register___U9354 ( .A1(register__n12282), .A2(register__n577), .B1(register__n10237), .B2(register__n590), 
        .Y(register__n13219) );
  INVx1_ASAP7_75t_R register___U9355 ( .A(register__n3659), .Y(register__n5942) );
  OA22x2_ASAP7_75t_R register___U9356 ( .A1(register__n12283), .A2(register__n103), .B1(register__n8732), .B2(register__n1142), 
        .Y(register__n13159) );
  INVx1_ASAP7_75t_R register___U9357 ( .A(register__n13159), .Y(register__n5943) );
  OA22x2_ASAP7_75t_R register___U9358 ( .A1(register__net63336), .A2(register__n1973), .B1(register__n10257), .B2(
        n11787), .Y(register__n12896) );
  INVx1_ASAP7_75t_R register___U9359 ( .A(register__n3330), .Y(register__n5945) );
  OA22x2_ASAP7_75t_R register___U9360 ( .A1(register__n12084), .A2(register__n118), .B1(register__n8833), .B2(register__n1194), 
        .Y(register__n13106) );
  INVx1_ASAP7_75t_R register___U9361 ( .A(register__n4088), .Y(register__n5946) );
  INVx3_ASAP7_75t_R register___U9362 ( .A(register__n12097), .Y(register__n12084) );
  OA22x2_ASAP7_75t_R register___U9363 ( .A1(register__net63264), .A2(register__n113), .B1(register__net90253), .B2(
        n1546), .Y(register__n12585) );
  INVx6_ASAP7_75t_R register___U9364 ( .A(register__net140283), .Y(register__net63264) );
  OA22x2_ASAP7_75t_R register___U9365 ( .A1(register__n12192), .A2(register__n11730), .B1(register__n10353), .B2(register__n1164), 
        .Y(register__n13373) );
  OA22x2_ASAP7_75t_R register___U9366 ( .A1(register__n12451), .A2(register__n3719), .B1(register__n9539), .B2(register__n1163), 
        .Y(register__n13359) );
  BUFx12f_ASAP7_75t_R register___U9367 ( .A(register__net64392), .Y(register__net64378) );
  OA22x2_ASAP7_75t_R register___U9368 ( .A1(register__n12032), .A2(register__n339), .B1(register__n9630), .B2(register__n344), 
        .Y(register__n12743) );
  INVx1_ASAP7_75t_R register___U9369 ( .A(register__n3575), .Y(register__n5949) );
  OA22x2_ASAP7_75t_R register___U9370 ( .A1(register__n3073), .A2(register__n1266), .B1(register__n9692), .B2(register__n3821), 
        .Y(register__n13144) );
  OA22x2_ASAP7_75t_R register___U9371 ( .A1(register__n5074), .A2(register__n702), .B1(register__n10347), .B2(register__n694), 
        .Y(register__n13327) );
  INVx1_ASAP7_75t_R register___U9372 ( .A(register__n4507), .Y(register__n5950) );
  INVx2_ASAP7_75t_R register___U9373 ( .A(register__n9373), .Y(register__n11437) );
  BUFx2_ASAP7_75t_R register___U9374 ( .A(register__C6422_net60224), .Y(register__net117114) );
  INVx2_ASAP7_75t_R register___U9375 ( .A(register__n8827), .Y(register__n11482) );
  BUFx2_ASAP7_75t_R register___U9376 ( .A(register__n10959), .Y(register__n5953) );
  BUFx2_ASAP7_75t_R register___U9377 ( .A(register__n10789), .Y(register__n5954) );
  BUFx2_ASAP7_75t_R register___U9378 ( .A(register__n11021), .Y(register__n5955) );
  INVx2_ASAP7_75t_R register___U9379 ( .A(register__n9559), .Y(register__n11108) );
  INVx2_ASAP7_75t_R register___U9380 ( .A(register__n9487), .Y(register__n10958) );
  INVx2_ASAP7_75t_R register___U9381 ( .A(register__n9493), .Y(register__n10870) );
  INVx2_ASAP7_75t_R register___U9382 ( .A(register__n9495), .Y(register__n10825) );
  INVx2_ASAP7_75t_R register___U9383 ( .A(register__n9499), .Y(register__n11204) );
  INVx2_ASAP7_75t_R register___U9384 ( .A(register__n9453), .Y(register__n10596) );
  INVx2_ASAP7_75t_R register___U9385 ( .A(register__n9571), .Y(register__n11455) );
  BUFx4f_ASAP7_75t_R register___U9386 ( .A(register__n9160), .Y(register__n5956) );
  BUFx6f_ASAP7_75t_R register___U9387 ( .A(register__n8688), .Y(register__n11306) );
  BUFx12f_ASAP7_75t_R register___U9388 ( .A(register__net112763), .Y(register__net116957) );
  INVx6_ASAP7_75t_R register___U9389 ( .A(register__n3387), .Y(register__n12080) );
  BUFx2_ASAP7_75t_R register___U9390 ( .A(register__n5959), .Y(register__n5958) );
  BUFx2_ASAP7_75t_R register___U9391 ( .A(register__n12560), .Y(register__n5959) );
  BUFx2_ASAP7_75t_R register___U9392 ( .A(register__n5961), .Y(register__n5960) );
  BUFx2_ASAP7_75t_R register___U9393 ( .A(register__n12576), .Y(register__n5961) );
  BUFx2_ASAP7_75t_R register___U9394 ( .A(register__n5963), .Y(register__n5962) );
  BUFx2_ASAP7_75t_R register___U9395 ( .A(register__n13007), .Y(register__n5963) );
  BUFx2_ASAP7_75t_R register___U9396 ( .A(register__n5965), .Y(register__n5964) );
  BUFx2_ASAP7_75t_R register___U9397 ( .A(register__n13298), .Y(register__n5965) );
  BUFx2_ASAP7_75t_R register___U9398 ( .A(register__n5967), .Y(register__n5966) );
  BUFx2_ASAP7_75t_R register___U9399 ( .A(register__n13302), .Y(register__n5967) );
  BUFx2_ASAP7_75t_R register___U9400 ( .A(register__n5971), .Y(register__n5970) );
  BUFx2_ASAP7_75t_R register___U9401 ( .A(register__n13205), .Y(register__n5971) );
  BUFx2_ASAP7_75t_R register___U9402 ( .A(register__n5973), .Y(register__n5972) );
  BUFx2_ASAP7_75t_R register___U9403 ( .A(register__n5975), .Y(register__n5974) );
  BUFx2_ASAP7_75t_R register___U9404 ( .A(register__n5978), .Y(register__n5977) );
  BUFx2_ASAP7_75t_R register___U9405 ( .A(register__n5980), .Y(register__n5979) );
  BUFx2_ASAP7_75t_R register___U9406 ( .A(register__n5982), .Y(register__n5981) );
  BUFx2_ASAP7_75t_R register___U9407 ( .A(register__n13289), .Y(register__n5982) );
  OR2x2_ASAP7_75t_R register___U9408 ( .A(register__n5984), .B(register__n5985), .Y(register__n5983) );
  BUFx2_ASAP7_75t_R register___U9409 ( .A(register__n6394), .Y(register__n5984) );
  OR2x2_ASAP7_75t_R register___U9410 ( .A(register__net64832), .B(register__n1990), .Y(register__n6395) );
  INVx1_ASAP7_75t_R register___U9411 ( .A(register__n3875), .Y(register__n5985) );
  NOR2x1p5_ASAP7_75t_R register___U9412 ( .A(register__net89713), .B(register__n11731), .Y(register__n6394) );
  OR2x2_ASAP7_75t_R register___U9413 ( .A(register__n5987), .B(register__n5988), .Y(register__n5986) );
  BUFx2_ASAP7_75t_R register___U9414 ( .A(register__n6397), .Y(register__n5987) );
  OR2x2_ASAP7_75t_R register___U9415 ( .A(register__net64414), .B(register__n3119), .Y(register__n6398) );
  INVx1_ASAP7_75t_R register___U9416 ( .A(register__n4192), .Y(register__n5988) );
  BUFx2_ASAP7_75t_R register___U9417 ( .A(register__n12988), .Y(register__n5989) );
  BUFx3_ASAP7_75t_R register___U9418 ( .A(register__n5991), .Y(register__n5990) );
  BUFx2_ASAP7_75t_R register___U9419 ( .A(register__n11543), .Y(register__n5991) );
  BUFx3_ASAP7_75t_R register___U9420 ( .A(register__n5993), .Y(register__n5992) );
  BUFx2_ASAP7_75t_R register___U9421 ( .A(register__n11546), .Y(register__n5993) );
  BUFx3_ASAP7_75t_R register___U9422 ( .A(register__n5997), .Y(register__n5996) );
  BUFx2_ASAP7_75t_R register___U9423 ( .A(register__n11244), .Y(register__n5997) );
  BUFx4f_ASAP7_75t_R register___U9424 ( .A(register__n11242), .Y(register__n7963) );
  INVx2_ASAP7_75t_R register___U9425 ( .A(register__n7963), .Y(register__n5998) );
  BUFx3_ASAP7_75t_R register___U9426 ( .A(register__n6002), .Y(register__n6001) );
  BUFx2_ASAP7_75t_R register___U9427 ( .A(register__n11159), .Y(register__n6002) );
  BUFx3_ASAP7_75t_R register___U9428 ( .A(register__n6004), .Y(register__n6003) );
  BUFx2_ASAP7_75t_R register___U9429 ( .A(register__n11157), .Y(register__n6004) );
  BUFx4f_ASAP7_75t_R register___U9430 ( .A(register__n6003), .Y(register__n9223) );
  BUFx3_ASAP7_75t_R register___U9431 ( .A(register__n6007), .Y(register__n6006) );
  BUFx2_ASAP7_75t_R register___U9432 ( .A(register__n11158), .Y(register__n6007) );
  BUFx3_ASAP7_75t_R register___U9433 ( .A(register__n11346), .Y(register__n6008) );
  BUFx3_ASAP7_75t_R register___U9434 ( .A(register__n6010), .Y(register__n6009) );
  BUFx2_ASAP7_75t_R register___U9435 ( .A(register__n11499), .Y(register__n6010) );
  BUFx3_ASAP7_75t_R register___U9436 ( .A(register__n6012), .Y(register__n6011) );
  BUFx2_ASAP7_75t_R register___U9437 ( .A(register__n11498), .Y(register__n6012) );
  INVx2_ASAP7_75t_R register___U9438 ( .A(register__n71), .Y(register__n6013) );
  BUFx3_ASAP7_75t_R register___U9439 ( .A(register__n6015), .Y(register__n6014) );
  BUFx2_ASAP7_75t_R register___U9440 ( .A(register__n11582), .Y(register__n6015) );
  BUFx3_ASAP7_75t_R register___U9441 ( .A(register__n6017), .Y(register__n6016) );
  BUFx2_ASAP7_75t_R register___U9442 ( .A(register__n11581), .Y(register__n6017) );
  BUFx4f_ASAP7_75t_R register___U9443 ( .A(register__n6018), .Y(register__n7972) );
  INVx2_ASAP7_75t_R register___U9444 ( .A(register__n7972), .Y(register__n6020) );
  BUFx3_ASAP7_75t_R register___U9445 ( .A(register__n6024), .Y(register__n6023) );
  BUFx2_ASAP7_75t_R register___U9446 ( .A(register__n11369), .Y(register__n6024) );
  BUFx2_ASAP7_75t_R register___U9447 ( .A(register__n9208), .Y(register__n6027) );
  BUFx3_ASAP7_75t_R register___U9448 ( .A(register__n6029), .Y(register__n6028) );
  BUFx3_ASAP7_75t_R register___U9449 ( .A(register__n6031), .Y(register__n6030) );
  BUFx2_ASAP7_75t_R register___U9450 ( .A(register__n11641), .Y(register__n6031) );
  BUFx4f_ASAP7_75t_R register___U9451 ( .A(register__n6030), .Y(register__n8327) );
  INVx2_ASAP7_75t_R register___U9452 ( .A(register__n8327), .Y(register__n6032) );
  OR2x2_ASAP7_75t_R register___U9453 ( .A(register__n6034), .B(register__n6035), .Y(register__n6033) );
  OR2x2_ASAP7_75t_R register___U9454 ( .A(register__net149934), .B(register__n11042), .Y(register__n8328) );
  INVx1_ASAP7_75t_R register___U9455 ( .A(register__n5117), .Y(register__n6034) );
  OR2x2_ASAP7_75t_R register___U9456 ( .A(register__n714), .B(register__n11645), .Y(register__n8329) );
  INVx1_ASAP7_75t_R register___U9457 ( .A(register__n5118), .Y(register__n6035) );
  BUFx3_ASAP7_75t_R register___U9458 ( .A(register__net91073), .Y(register__net116359) );
  BUFx4f_ASAP7_75t_R register___U9459 ( .A(register__net91073), .Y(register__net116361) );
  BUFx3_ASAP7_75t_R register___U9460 ( .A(register__n6843), .Y(register__n6036) );
  BUFx3_ASAP7_75t_R register___U9461 ( .A(register__n6540), .Y(register__n6037) );
  BUFx3_ASAP7_75t_R register___U9462 ( .A(register__n10014), .Y(register__n6038) );
  BUFx4f_ASAP7_75t_R register___U9463 ( .A(register__n10014), .Y(register__n6039) );
  BUFx2_ASAP7_75t_R register___U9464 ( .A(register__n10014), .Y(register__n6040) );
  BUFx3_ASAP7_75t_R register___U9465 ( .A(register__n8122), .Y(register__n6041) );
  BUFx6f_ASAP7_75t_R register___U9466 ( .A(register__n8121), .Y(register__n10152) );
  BUFx4f_ASAP7_75t_R register___U9467 ( .A(register__n6041), .Y(register__n8121) );
  BUFx3_ASAP7_75t_R register___U9468 ( .A(register__n6545), .Y(register__n6042) );
  BUFx3_ASAP7_75t_R register___U9469 ( .A(register__n8148), .Y(register__n6043) );
  BUFx6f_ASAP7_75t_R register___U9470 ( .A(register__n8147), .Y(register__n10218) );
  BUFx4f_ASAP7_75t_R register___U9471 ( .A(register__n6043), .Y(register__n8147) );
  BUFx12f_ASAP7_75t_R register___U9472 ( .A(register__n9811), .Y(register__n6045) );
  BUFx6f_ASAP7_75t_R register___U9473 ( .A(register__n10506), .Y(register__n10505) );
  BUFx3_ASAP7_75t_R register___U9474 ( .A(register__n7209), .Y(register__n6046) );
  BUFx12f_ASAP7_75t_R register___U9475 ( .A(register__net64728), .Y(register__net64708) );
  BUFx2_ASAP7_75t_R register___U9476 ( .A(Reg_data[612]), .Y(register__n6047) );
  BUFx6f_ASAP7_75t_R register___U9477 ( .A(register__n9962), .Y(register__n9961) );
  BUFx4f_ASAP7_75t_R register___U9478 ( .A(register__n5646), .Y(register__n9962) );
  BUFx2_ASAP7_75t_R register___U9479 ( .A(Reg_data[528]), .Y(register__n6048) );
  BUFx6f_ASAP7_75t_R register___U9480 ( .A(register__n9424), .Y(register__n9423) );
  BUFx4f_ASAP7_75t_R register___U9481 ( .A(register__n5647), .Y(register__n9424) );
  BUFx2_ASAP7_75t_R register___U9482 ( .A(Reg_data[163]), .Y(register__n6049) );
  BUFx4f_ASAP7_75t_R register___U9483 ( .A(register__n10012), .Y(register__n6050) );
  BUFx2_ASAP7_75t_R register___U9484 ( .A(register__n10012), .Y(register__n6051) );
  BUFx6f_ASAP7_75t_R register___U9485 ( .A(register__n10013), .Y(register__n10012) );
  BUFx4f_ASAP7_75t_R register___U9486 ( .A(register__n5651), .Y(register__n10013) );
  BUFx2_ASAP7_75t_R register___U9487 ( .A(Reg_data[393]), .Y(register__n6052) );
  BUFx6f_ASAP7_75t_R register___U9488 ( .A(register__n10435), .Y(register__n10434) );
  BUFx4f_ASAP7_75t_R register___U9489 ( .A(register__n5510), .Y(register__n10435) );
  BUFx2_ASAP7_75t_R register___U9490 ( .A(Reg_data[51]), .Y(register__n6053) );
  BUFx6f_ASAP7_75t_R register___U9491 ( .A(register__n10159), .Y(register__n10158) );
  BUFx4f_ASAP7_75t_R register___U9492 ( .A(register__n5832), .Y(register__n10159) );
  BUFx2_ASAP7_75t_R register___U9493 ( .A(Reg_data[524]), .Y(register__n6054) );
  BUFx6f_ASAP7_75t_R register___U9494 ( .A(register__n9434), .Y(register__n9433) );
  BUFx4f_ASAP7_75t_R register___U9495 ( .A(register__n5512), .Y(register__n9434) );
  BUFx2_ASAP7_75t_R register___U9496 ( .A(Reg_data[443]), .Y(register__n6055) );
  BUFx6f_ASAP7_75t_R register___U9497 ( .A(register__n10443), .Y(register__n10442) );
  BUFx4f_ASAP7_75t_R register___U9498 ( .A(register__n5837), .Y(register__n10443) );
  INVx1_ASAP7_75t_R register___U9499 ( .A(register__n5737), .Y(register__n6056) );
  INVx1_ASAP7_75t_R register___U9500 ( .A(register__n5745), .Y(register__n6058) );
  BUFx3_ASAP7_75t_R register___U9501 ( .A(register__net116147), .Y(register__net116146) );
  BUFx2_ASAP7_75t_R register___U9502 ( .A(Reg_data[985]), .Y(register__net116147) );
  BUFx3_ASAP7_75t_R register___U9503 ( .A(register__net116143), .Y(register__net116142) );
  BUFx2_ASAP7_75t_R register___U9504 ( .A(Reg_data[965]), .Y(register__net116143) );
  BUFx3_ASAP7_75t_R register___U9505 ( .A(register__n6061), .Y(register__n6060) );
  BUFx2_ASAP7_75t_R register___U9506 ( .A(Reg_data[962]), .Y(register__n6061) );
  BUFx3_ASAP7_75t_R register___U9507 ( .A(register__n6063), .Y(register__n6062) );
  BUFx2_ASAP7_75t_R register___U9508 ( .A(Reg_data[960]), .Y(register__n6063) );
  BUFx3_ASAP7_75t_R register___U9509 ( .A(register__n6065), .Y(register__n6064) );
  BUFx2_ASAP7_75t_R register___U9510 ( .A(Reg_data[932]), .Y(register__n6065) );
  BUFx3_ASAP7_75t_R register___U9511 ( .A(register__n6067), .Y(register__n6066) );
  BUFx2_ASAP7_75t_R register___U9512 ( .A(Reg_data[928]), .Y(register__n6067) );
  BUFx3_ASAP7_75t_R register___U9513 ( .A(register__n6069), .Y(register__n6068) );
  BUFx2_ASAP7_75t_R register___U9514 ( .A(Reg_data[904]), .Y(register__n6069) );
  BUFx3_ASAP7_75t_R register___U9515 ( .A(register__n6071), .Y(register__n6070) );
  BUFx2_ASAP7_75t_R register___U9516 ( .A(Reg_data[900]), .Y(register__n6071) );
  BUFx3_ASAP7_75t_R register___U9517 ( .A(register__n6073), .Y(register__n6072) );
  BUFx2_ASAP7_75t_R register___U9518 ( .A(Reg_data[816]), .Y(register__n6073) );
  BUFx3_ASAP7_75t_R register___U9519 ( .A(register__net116111), .Y(register__net116110) );
  BUFx2_ASAP7_75t_R register___U9520 ( .A(Reg_data[806]), .Y(register__net116111) );
  BUFx3_ASAP7_75t_R register___U9521 ( .A(register__n6075), .Y(register__n6074) );
  BUFx2_ASAP7_75t_R register___U9522 ( .A(Reg_data[803]), .Y(register__n6075) );
  BUFx3_ASAP7_75t_R register___U9523 ( .A(register__n6077), .Y(register__n6076) );
  BUFx2_ASAP7_75t_R register___U9524 ( .A(Reg_data[802]), .Y(register__n6077) );
  BUFx3_ASAP7_75t_R register___U9525 ( .A(register__n6079), .Y(register__n6078) );
  BUFx2_ASAP7_75t_R register___U9526 ( .A(Reg_data[800]), .Y(register__n6079) );
  BUFx3_ASAP7_75t_R register___U9527 ( .A(register__n6081), .Y(register__n6080) );
  BUFx2_ASAP7_75t_R register___U9528 ( .A(Reg_data[726]), .Y(register__n6081) );
  BUFx3_ASAP7_75t_R register___U9529 ( .A(register__n6083), .Y(register__n6082) );
  BUFx2_ASAP7_75t_R register___U9530 ( .A(Reg_data[693]), .Y(register__n6083) );
  BUFx3_ASAP7_75t_R register___U9531 ( .A(register__n6085), .Y(register__n6084) );
  BUFx2_ASAP7_75t_R register___U9532 ( .A(Reg_data[641]), .Y(register__n6085) );
  BUFx3_ASAP7_75t_R register___U9533 ( .A(register__n6087), .Y(register__n6086) );
  BUFx2_ASAP7_75t_R register___U9534 ( .A(Reg_data[534]), .Y(register__n6087) );
  BUFx3_ASAP7_75t_R register___U9535 ( .A(register__n6089), .Y(register__n6088) );
  BUFx2_ASAP7_75t_R register___U9536 ( .A(Reg_data[469]), .Y(register__n6089) );
  BUFx3_ASAP7_75t_R register___U9537 ( .A(register__net116075), .Y(register__net116074) );
  BUFx2_ASAP7_75t_R register___U9538 ( .A(Reg_data[454]), .Y(register__net116075) );
  BUFx3_ASAP7_75t_R register___U9539 ( .A(register__n6091), .Y(register__n6090) );
  BUFx2_ASAP7_75t_R register___U9540 ( .A(Reg_data[452]), .Y(register__n6091) );
  BUFx3_ASAP7_75t_R register___U9541 ( .A(register__n6093), .Y(register__n6092) );
  BUFx2_ASAP7_75t_R register___U9542 ( .A(Reg_data[210]), .Y(register__n6093) );
  BUFx3_ASAP7_75t_R register___U9543 ( .A(register__n6095), .Y(register__n6094) );
  BUFx2_ASAP7_75t_R register___U9544 ( .A(Reg_data[973]), .Y(register__n6095) );
  BUFx3_ASAP7_75t_R register___U9545 ( .A(register__n9264), .Y(register__n6096) );
  BUFx2_ASAP7_75t_R register___U9546 ( .A(register__n9264), .Y(register__n6097) );
  BUFx4f_ASAP7_75t_R register___U9547 ( .A(register__n9264), .Y(register__n6098) );
  BUFx3_ASAP7_75t_R register___U9548 ( .A(register__n6100), .Y(register__n6099) );
  BUFx2_ASAP7_75t_R register___U9549 ( .A(Reg_data[828]), .Y(register__n6100) );
  BUFx3_ASAP7_75t_R register___U9550 ( .A(register__n6102), .Y(register__n6101) );
  BUFx2_ASAP7_75t_R register___U9551 ( .A(Reg_data[991]), .Y(register__n6102) );
  BUFx3_ASAP7_75t_R register___U9552 ( .A(register__net116045), .Y(register__net116044) );
  BUFx2_ASAP7_75t_R register___U9553 ( .A(Reg_data[984]), .Y(register__net116045) );
  BUFx3_ASAP7_75t_R register___U9554 ( .A(register__net116041), .Y(register__net116040) );
  BUFx2_ASAP7_75t_R register___U9555 ( .A(Reg_data[975]), .Y(register__net116041) );
  BUFx3_ASAP7_75t_R register___U9556 ( .A(register__n6104), .Y(register__n6103) );
  BUFx2_ASAP7_75t_R register___U9557 ( .A(Reg_data[827]), .Y(register__n6104) );
  BUFx3_ASAP7_75t_R register___U9558 ( .A(register__n6106), .Y(register__n6105) );
  BUFx2_ASAP7_75t_R register___U9559 ( .A(Reg_data[974]), .Y(register__n6106) );
  BUFx3_ASAP7_75t_R register___U9560 ( .A(register__n6108), .Y(register__n6107) );
  BUFx2_ASAP7_75t_R register___U9561 ( .A(Reg_data[703]), .Y(register__n6108) );
  BUFx3_ASAP7_75t_R register___U9562 ( .A(register__net116025), .Y(register__net116024) );
  BUFx2_ASAP7_75t_R register___U9563 ( .A(Reg_data[317]), .Y(register__net116025) );
  BUFx3_ASAP7_75t_R register___U9564 ( .A(register__n6110), .Y(register__n6109) );
  BUFx2_ASAP7_75t_R register___U9565 ( .A(Reg_data[717]), .Y(register__n6110) );
  BUFx3_ASAP7_75t_R register___U9566 ( .A(register__n10134), .Y(register__n6111) );
  BUFx2_ASAP7_75t_R register___U9567 ( .A(register__n10134), .Y(register__n6112) );
  BUFx4f_ASAP7_75t_R register___U9568 ( .A(register__n10134), .Y(register__n6113) );
  BUFx3_ASAP7_75t_R register___U9569 ( .A(register__n6115), .Y(register__n6114) );
  BUFx2_ASAP7_75t_R register___U9570 ( .A(Reg_data[199]), .Y(register__n6115) );
  BUFx3_ASAP7_75t_R register___U9571 ( .A(register__n6117), .Y(register__n6116) );
  BUFx2_ASAP7_75t_R register___U9572 ( .A(Reg_data[7]), .Y(register__n6117) );
  BUFx3_ASAP7_75t_R register___U9573 ( .A(register__net115997), .Y(register__net115996) );
  BUFx2_ASAP7_75t_R register___U9574 ( .A(Reg_data[719]), .Y(register__net115997) );
  BUFx2_ASAP7_75t_R register___U9575 ( .A(register__net89393), .Y(register__net115999) );
  BUFx4f_ASAP7_75t_R register___U9576 ( .A(register__net89393), .Y(register__net116000) );
  BUFx3_ASAP7_75t_R register___U9577 ( .A(register__net115993), .Y(register__net115992) );
  BUFx2_ASAP7_75t_R register___U9578 ( .A(Reg_data[431]), .Y(register__net115993) );
  BUFx3_ASAP7_75t_R register___U9579 ( .A(register__n6119), .Y(register__n6118) );
  BUFx2_ASAP7_75t_R register___U9580 ( .A(Reg_data[574]), .Y(register__n6119) );
  BUFx3_ASAP7_75t_R register___U9581 ( .A(register__net115985), .Y(register__net115984) );
  BUFx2_ASAP7_75t_R register___U9582 ( .A(Reg_data[682]), .Y(register__net115985) );
  BUFx3_ASAP7_75t_R register___U9583 ( .A(register__net115975), .Y(register__net115974) );
  BUFx2_ASAP7_75t_R register___U9584 ( .A(Reg_data[714]), .Y(register__net115975) );
  BUFx2_ASAP7_75t_R register___U9585 ( .A(register__net89273), .Y(register__net115976) );
  BUFx4f_ASAP7_75t_R register___U9586 ( .A(register__net89273), .Y(register__net115978) );
  BUFx3_ASAP7_75t_R register___U9587 ( .A(register__n6121), .Y(register__n6120) );
  BUFx2_ASAP7_75t_R register___U9588 ( .A(Reg_data[727]), .Y(register__n6121) );
  BUFx3_ASAP7_75t_R register___U9589 ( .A(register__n6123), .Y(register__n6122) );
  BUFx2_ASAP7_75t_R register___U9590 ( .A(Reg_data[471]), .Y(register__n6123) );
  BUFx3_ASAP7_75t_R register___U9591 ( .A(register__n6125), .Y(register__n6124) );
  BUFx2_ASAP7_75t_R register___U9592 ( .A(Reg_data[831]), .Y(register__n6125) );
  BUFx12f_ASAP7_75t_R register___U9593 ( .A(register__net121483), .Y(register__net62858) );
  INVx2_ASAP7_75t_R register___U9594 ( .A(register__n12468), .Y(register__n12452) );
  BUFx6f_ASAP7_75t_R register___U9595 ( .A(register__n5224), .Y(register__n12468) );
  BUFx12f_ASAP7_75t_R register___U9596 ( .A(register__n3448), .Y(register__n12473) );
  OA22x2_ASAP7_75t_R register___U9597 ( .A1(register__n12053), .A2(register__n986), .B1(register__n10090), .B2(register__n975), 
        .Y(register__n13200) );
  OA22x2_ASAP7_75t_R register___U9598 ( .A1(register__net129768), .A2(register__n701), .B1(register__n9513), .B2(register__n671), 
        .Y(register__n13328) );
  OA22x2_ASAP7_75t_R register___U9599 ( .A1(register__net64348), .A2(register__n1003), .B1(register__net89581), .B2(
        n975), .Y(register__n13197) );
  INVx1_ASAP7_75t_R register___U9600 ( .A(register__n4009), .Y(register__n6128) );
  OA22x2_ASAP7_75t_R register___U9601 ( .A1(register__net63238), .A2(register__n700), .B1(register__net91331), .B2(register__n686), .Y(register__n13313) );
  INVx3_ASAP7_75t_R register___U9602 ( .A(register__net63272), .Y(register__net63238) );
  OA22x2_ASAP7_75t_R register___U9603 ( .A1(register__n12080), .A2(register__n1988), .B1(register__n10273), .B2(register__n4952), 
        .Y(register__n13352) );
  OA22x2_ASAP7_75t_R register___U9604 ( .A1(register__n12082), .A2(register__n577), .B1(register__n8351), .B2(register__n584), 
        .Y(register__n13229) );
  OA22x2_ASAP7_75t_R register___U9605 ( .A1(register__n12170), .A2(register__n955), .B1(register__n9907), .B2(register__n959), 
        .Y(register__n13025) );
  OA22x2_ASAP7_75t_R register___U9606 ( .A1(register__n12310), .A2(register__n1989), .B1(register__n10078), .B2(register__n4374), 
        .Y(register__n13343) );
  OA22x2_ASAP7_75t_R register___U9607 ( .A1(register__n12145), .A2(register__n575), .B1(register__n10124), .B2(register__n580), 
        .Y(register__n13225) );
  INVx6_ASAP7_75t_R register___U9608 ( .A(register__n12156), .Y(register__n12145) );
  OA22x2_ASAP7_75t_R register___U9609 ( .A1(register__n12404), .A2(register__n1794), .B1(register__n10291), .B2(register__n1630), 
        .Y(register__n12751) );
  INVx1_ASAP7_75t_R register___U9610 ( .A(register__n5095), .Y(register__n6131) );
  OA22x2_ASAP7_75t_R register___U9611 ( .A1(register__n12234), .A2(register__n1792), .B1(register__n10317), .B2(register__n1633), 
        .Y(register__n12760) );
  OA22x2_ASAP7_75t_R register___U9612 ( .A1(register__n12339), .A2(register__n575), .B1(register__n7459), .B2(register__n579), 
        .Y(register__n13217) );
  INVx1_ASAP7_75t_R register___U9613 ( .A(register__n5570), .Y(register__n6133) );
  OA22x2_ASAP7_75t_R register___U9614 ( .A1(register__n11983), .A2(register__n1989), .B1(register__n8945), .B2(register__n5183), 
        .Y(register__n13355) );
  OA22x2_ASAP7_75t_R register___U9615 ( .A1(register__net62664), .A2(register__n460), .B1(register__n6377), .B2(register__n469), 
        .Y(register__n12919) );
  INVx6_ASAP7_75t_R register___U9616 ( .A(register__net63274), .Y(register__net63242) );
  OA22x2_ASAP7_75t_R register___U9617 ( .A1(register__net64418), .A2(register__n575), .B1(register__net103455), .B2(
        n588), .Y(register__n13228) );
  OA22x2_ASAP7_75t_R register___U9618 ( .A1(register__net63336), .A2(register__n460), .B1(register__n7217), .B2(register__n466), 
        .Y(register__n12926) );
  INVx1_ASAP7_75t_R register___U9619 ( .A(register__n4783), .Y(register__n6137) );
  OA22x2_ASAP7_75t_R register___U9620 ( .A1(register__n12090), .A2(register__n1794), .B1(register__n8522), .B2(register__n1641), 
        .Y(register__n12767) );
  INVx1_ASAP7_75t_R register___U9621 ( .A(register__n12767), .Y(register__n6138) );
  OA22x2_ASAP7_75t_R register___U9622 ( .A1(register__net64350), .A2(register__n1647), .B1(register__net89593), .B2(
        n1632), .Y(register__n12765) );
  OA22x2_ASAP7_75t_R register___U9623 ( .A1(register__n12454), .A2(register__n576), .B1(register__n10191), .B2(register__n584), 
        .Y(register__n13209) );
  INVx4_ASAP7_75t_R register___U9624 ( .A(register__n12469), .Y(register__n12454) );
  BUFx12f_ASAP7_75t_R register___U9625 ( .A(register__n11806), .Y(register__n11891) );
  INVx1_ASAP7_75t_R register___U9626 ( .A(register__n4340), .Y(register__n6141) );
  AND4x1_ASAP7_75t_R register___U9627 ( .A(register__n6140), .B(register__n6827), .C(register__n4338), .D(register__n6141), .Y(
        n10634) );
  INVx1_ASAP7_75t_R register___U9628 ( .A(register__n4361), .Y(register__n6143) );
  INVx1_ASAP7_75t_R register___U9629 ( .A(register__n4363), .Y(register__n6144) );
  INVx1_ASAP7_75t_R register___U9630 ( .A(register__n4365), .Y(register__n6145) );
  INVx1_ASAP7_75t_R register___U9631 ( .A(register__n5411), .Y(register__n6146) );
  INVx1_ASAP7_75t_R register___U9632 ( .A(register__n10943), .Y(register__n6147) );
  INVx1_ASAP7_75t_R register___U9633 ( .A(register__n10945), .Y(register__n6148) );
  INVx1_ASAP7_75t_R register___U9634 ( .A(register__n3985), .Y(register__n6149) );
  INVx1_ASAP7_75t_R register___U9635 ( .A(register__n4460), .Y(register__n6150) );
  INVx1_ASAP7_75t_R register___U9636 ( .A(register__n4464), .Y(register__n6152) );
  INVx1_ASAP7_75t_R register___U9637 ( .A(register__n4456), .Y(register__n6153) );
  INVx1_ASAP7_75t_R register___U9638 ( .A(register__n4458), .Y(register__n6154) );
  AND4x1_ASAP7_75t_R register___U9639 ( .A(register__n6154), .B(register__n1614), .C(register__n1804), .D(register__n4457), .Y(
        n10733) );
  INVx1_ASAP7_75t_R register___U9640 ( .A(register__n5423), .Y(register__n6155) );
  INVx1_ASAP7_75t_R register___U9641 ( .A(register__n5425), .Y(register__n6156) );
  INVx1_ASAP7_75t_R register___U9642 ( .A(register__n5427), .Y(register__n6157) );
  INVx1_ASAP7_75t_R register___U9643 ( .A(register__n4560), .Y(register__n6158) );
  INVx1_ASAP7_75t_R register___U9644 ( .A(register__n4563), .Y(register__n6159) );
  OA22x2_ASAP7_75t_R register___U9645 ( .A1(register__n12255), .A2(register__n1416), .B1(register__n7436), .B2(register__n1419), 
        .Y(register__n12992) );
  INVx1_ASAP7_75t_R register___U9646 ( .A(register__n4132), .Y(register__n6163) );
  OA22x2_ASAP7_75t_R register___U9647 ( .A1(register__n12366), .A2(register__n399), .B1(register__n8029), .B2(register__n3416), 
        .Y(register__n13294) );
  INVx1_ASAP7_75t_R register___U9648 ( .A(register__n4655), .Y(register__n6164) );
  OA22x2_ASAP7_75t_R register___U9649 ( .A1(register__net62990), .A2(register__n578), .B1(register__n8200), .B2(register__n582), 
        .Y(register__n13212) );
  OA22x2_ASAP7_75t_R register___U9650 ( .A1(register__n12057), .A2(register__n462), .B1(register__n7994), .B2(register__n465), 
        .Y(register__n12941) );
  OA22x2_ASAP7_75t_R register___U9651 ( .A1(register__n12263), .A2(register__n4033), .B1(register__n8805), .B2(register__n11841), 
        .Y(register__n12535) );
  INVx1_ASAP7_75t_R register___U9652 ( .A(register__n5403), .Y(register__n6165) );
  OA22x2_ASAP7_75t_R register___U9653 ( .A1(register__n12317), .A2(register__n1413), .B1(register__n7988), .B2(register__n1419), 
        .Y(register__n12990) );
  INVx1_ASAP7_75t_R register___U9654 ( .A(register__n5268), .Y(register__n6166) );
  OA22x2_ASAP7_75t_R register___U9655 ( .A1(register__n12378), .A2(register__n4033), .B1(register__n9248), .B2(register__n11843), 
        .Y(register__n12531) );
  INVx1_ASAP7_75t_R register___U9656 ( .A(register__n5564), .Y(register__n6168) );
  OA22x2_ASAP7_75t_R register___U9657 ( .A1(register__n11964), .A2(register__n4033), .B1(register__n9329), .B2(register__n4844), 
        .Y(register__n12551) );
  OA22x2_ASAP7_75t_R register___U9658 ( .A1(register__n12261), .A2(register__n116), .B1(register__n7984), .B2(register__n1673), 
        .Y(register__n12645) );
  INVx1_ASAP7_75t_R register___U9659 ( .A(register__n3712), .Y(register__n6170) );
  OA22x2_ASAP7_75t_R register___U9660 ( .A1(register__n12320), .A2(register__n1647), .B1(register__n9919), .B2(register__n1617), 
        .Y(register__n12757) );
  INVx1_ASAP7_75t_R register___U9661 ( .A(register__n5075), .Y(register__n6171) );
  OA22x2_ASAP7_75t_R register___U9662 ( .A1(register__n12259), .A2(register__n1647), .B1(register__n9921), .B2(register__n1637), 
        .Y(register__n12759) );
  INVx1_ASAP7_75t_R register___U9663 ( .A(register__n3884), .Y(register__n6172) );
  OA22x2_ASAP7_75t_R register___U9664 ( .A1(register__net64770), .A2(register__n1794), .B1(register__net90149), .B2(
        n1636), .Y(register__n12770) );
  OA22x2_ASAP7_75t_R register___U9665 ( .A1(register__net64854), .A2(register__n1793), .B1(register__net90145), .B2(
        n1621), .Y(register__n12771) );
  OA22x2_ASAP7_75t_R register___U9666 ( .A1(register__n11994), .A2(register__n104), .B1(register__n9925), .B2(register__n1619), 
        .Y(register__n12774) );
  OA22x2_ASAP7_75t_R register___U9667 ( .A1(register__n11931), .A2(register__n1647), .B1(register__n9927), .B2(register__n1635), 
        .Y(register__n12776) );
  INVx1_ASAP7_75t_R register___U9668 ( .A(register__n4130), .Y(register__n6177) );
  OA22x2_ASAP7_75t_R register___U9669 ( .A1(register__net63168), .A2(register__n459), .B1(register__net89969), .B2(register__n464), .Y(register__n12924) );
  OA22x2_ASAP7_75t_R register___U9670 ( .A1(register__net64848), .A2(register__n459), .B1(register__net89953), .B2(register__n468), .Y(register__n12944) );
  OA22x2_ASAP7_75t_R register___U9671 ( .A1(register__net64920), .A2(register__n459), .B1(register__n9993), .B2(register__n464), 
        .Y(register__n12945) );
  INVx1_ASAP7_75t_R register___U9672 ( .A(register__n5751), .Y(register__n6178) );
  OA22x2_ASAP7_75t_R register___U9673 ( .A1(register__n11991), .A2(register__n461), .B1(register__n9425), .B2(register__n468), 
        .Y(register__n12947) );
  INVx1_ASAP7_75t_R register___U9674 ( .A(register__n4777), .Y(register__n6179) );
  OA22x2_ASAP7_75t_R register___U9675 ( .A1(register__n11957), .A2(register__n461), .B1(register__n10450), .B2(register__n463), 
        .Y(register__n12948) );
  OA22x2_ASAP7_75t_R register___U9676 ( .A1(register__net142928), .A2(register__n1416), .B1(register__net96895), .B2(
        n1419), .Y(register__n13004) );
  OA22x2_ASAP7_75t_R register___U9677 ( .A1(register__n11985), .A2(register__n2851), .B1(register__n10028), .B2(register__n3296), 
        .Y(register__n13283) );
  OA22x2_ASAP7_75t_R register___U9678 ( .A1(register__n12367), .A2(register__n577), .B1(register__n10052), .B2(register__n581), 
        .Y(register__n13216) );
  INVx1_ASAP7_75t_R register___U9679 ( .A(register__n4136), .Y(register__n6181) );
  OA22x2_ASAP7_75t_R register___U9680 ( .A1(register__n11924), .A2(register__n578), .B1(register__n10062), .B2(register__n590), 
        .Y(register__n13238) );
  OA22x2_ASAP7_75t_R register___U9681 ( .A1(register__n3700), .A2(register__n576), .B1(register__n9431), .B2(register__n585), .Y(
        n13236) );
  INVx1_ASAP7_75t_R register___U9682 ( .A(register__n4519), .Y(register__n6183) );
  OA22x2_ASAP7_75t_R register___U9683 ( .A1(register__net63338), .A2(register__n2823), .B1(register__n8724), .B2(register__n1926), 
        .Y(register__n12866) );
  OA22x2_ASAP7_75t_R register___U9684 ( .A1(register__net63000), .A2(register__n459), .B1(register__n8819), .B2(register__n470), 
        .Y(register__n12923) );
  OA22x2_ASAP7_75t_R register___U9685 ( .A1(register__n12226), .A2(register__n700), .B1(register__n10381), .B2(register__n695), 
        .Y(register__n13319) );
  OA22x2_ASAP7_75t_R register___U9686 ( .A1(register__n12168), .A2(register__n576), .B1(register__n10193), .B2(register__n582), 
        .Y(register__n13224) );
  OA22x2_ASAP7_75t_R register___U9687 ( .A1(register__n12280), .A2(register__n700), .B1(register__n10397), .B2(register__n687), 
        .Y(register__n13317) );
  INVx1_ASAP7_75t_R register___U9688 ( .A(register__n5011), .Y(register__n6186) );
  OA22x2_ASAP7_75t_R register___U9689 ( .A1(register__n12083), .A2(register__n1137), .B1(register__n8736), .B2(register__n1058), 
        .Y(register__n13167) );
  OA22x2_ASAP7_75t_R register___U9690 ( .A1(register__n12405), .A2(register__n3022), .B1(register__n7334), .B2(register__n1588), 
        .Y(register__n12695) );
  INVx1_ASAP7_75t_R register___U9691 ( .A(register__n5789), .Y(register__n6189) );
  OA22x2_ASAP7_75t_R register___U9692 ( .A1(register__n12395), .A2(register__n702), .B1(register__n10407), .B2(register__n670), 
        .Y(register__n13311) );
  OA22x2_ASAP7_75t_R register___U9693 ( .A1(register__net62662), .A2(register__n1416), .B1(register__n7390), .B2(register__n1417), 
        .Y(register__n12980) );
  INVx1_ASAP7_75t_R register___U9694 ( .A(register__n3033), .Y(register__n6191) );
  INVx1_ASAP7_75t_R register___U9695 ( .A(register__n3035), .Y(register__n6192) );
  INVx1_ASAP7_75t_R register___U9696 ( .A(register__n3008), .Y(register__n6194) );
  INVx1_ASAP7_75t_R register___U9697 ( .A(register__n3131), .Y(register__n6199) );
  OA22x2_ASAP7_75t_R register___U9698 ( .A1(register__net147310), .A2(register__n460), .B1(register__net91563), .B2(
        n465), .Y(register__n12943) );
  INVx1_ASAP7_75t_R register___U9699 ( .A(register__n3949), .Y(register__n6200) );
  OA22x2_ASAP7_75t_R register___U9700 ( .A1(register__n12368), .A2(register__n1568), .B1(register__n8825), .B2(register__n1198), 
        .Y(register__n13093) );
  INVx1_ASAP7_75t_R register___U9701 ( .A(register__n3767), .Y(register__n6201) );
  OA22x2_ASAP7_75t_R register___U9702 ( .A1(register__n3666), .A2(register__n1755), .B1(register__n9694), .B2(register__n3821), 
        .Y(register__n13145) );
  INVx1_ASAP7_75t_R register___U9703 ( .A(register__n2941), .Y(register__n6202) );
  OA22x2_ASAP7_75t_R register___U9704 ( .A1(register__n4864), .A2(register__n700), .B1(register__n9491), .B2(register__n680), .Y(
        n13316) );
  INVx2_ASAP7_75t_R register___U9705 ( .A(register__n12325), .Y(register__n12311) );
  OA22x2_ASAP7_75t_R register___U9706 ( .A1(register__n12019), .A2(register__n698), .B1(register__n9497), .B2(register__n689), 
        .Y(register__n13332) );
  INVx1_ASAP7_75t_R register___U9707 ( .A(register__n3928), .Y(register__n6204) );
  BUFx2_ASAP7_75t_R register___U9708 ( .A(register__n11482), .Y(register__n6205) );
  BUFx2_ASAP7_75t_R register___U9709 ( .A(register__n11437), .Y(register__n6206) );
  INVx2_ASAP7_75t_R register___U9710 ( .A(register__n9439), .Y(register__n10664) );
  BUFx2_ASAP7_75t_R register___U9711 ( .A(register__n11247), .Y(register__n6207) );
  BUFx2_ASAP7_75t_R register___U9712 ( .A(register__n11183), .Y(register__n6209) );
  BUFx2_ASAP7_75t_R register___U9713 ( .A(register__n10600), .Y(register__n6210) );
  INVx2_ASAP7_75t_R register___U9714 ( .A(register__n10377), .Y(register__n10766) );
  BUFx2_ASAP7_75t_R register___U9715 ( .A(register__n11108), .Y(register__n6211) );
  BUFx2_ASAP7_75t_R register___U9716 ( .A(register__n11353), .Y(register__n6213) );
  INVx2_ASAP7_75t_R register___U9717 ( .A(register__n10375), .Y(register__n11065) );
  INVx2_ASAP7_75t_R register___U9718 ( .A(register__n8829), .Y(register__n11415) );
  BUFx2_ASAP7_75t_R register___U9719 ( .A(register__n10825), .Y(register__n6215) );
  BUFx2_ASAP7_75t_R register___U9720 ( .A(register__n10870), .Y(register__n6216) );
  BUFx2_ASAP7_75t_R register___U9721 ( .A(register__n10958), .Y(register__n6218) );
  BUFx2_ASAP7_75t_R register___U9722 ( .A(register__n10764), .Y(register__n6220) );
  BUFx2_ASAP7_75t_R register___U9723 ( .A(register__C6422_net59833), .Y(register__net115136) );
  BUFx2_ASAP7_75t_R register___U9724 ( .A(register__n10846), .Y(register__n6221) );
  BUFx2_ASAP7_75t_R register___U9725 ( .A(register__n10684), .Y(register__n6222) );
  BUFx2_ASAP7_75t_R register___U9726 ( .A(register__n10892), .Y(register__n6223) );
  BUFx2_ASAP7_75t_R register___U9727 ( .A(register__n10742), .Y(register__n6224) );
  BUFx2_ASAP7_75t_R register___U9728 ( .A(register__n11414), .Y(register__n6225) );
  BUFx2_ASAP7_75t_R register___U9729 ( .A(register__n11020), .Y(register__n6226) );
  INVx2_ASAP7_75t_R register___U9730 ( .A(register__n9555), .Y(register__n11106) );
  BUFx2_ASAP7_75t_R register___U9731 ( .A(register__n11566), .Y(register__n6227) );
  BUFx2_ASAP7_75t_R register___U9732 ( .A(register__n10530), .Y(register__n6228) );
  INVx2_ASAP7_75t_R register___U9733 ( .A(register__n9451), .Y(register__n11327) );
  BUFx2_ASAP7_75t_R register___U9734 ( .A(register__n10935), .Y(register__n6229) );
  BUFx2_ASAP7_75t_R register___U9735 ( .A(register__n10914), .Y(register__n6230) );
  INVx2_ASAP7_75t_R register___U9736 ( .A(register__n9455), .Y(register__n11202) );
  BUFx2_ASAP7_75t_R register___U9737 ( .A(register__n11455), .Y(register__n6231) );
  BUFx2_ASAP7_75t_R register___U9738 ( .A(register__n11622), .Y(register__n6232) );
  INVx2_ASAP7_75t_R register___U9739 ( .A(register__n9529), .Y(register__n10741) );
  BUFx4f_ASAP7_75t_R register___U9740 ( .A(register__n10980), .Y(register__n6233) );
  BUFx2_ASAP7_75t_R register___U9741 ( .A(register__n8571), .Y(register__n6234) );
  BUFx3_ASAP7_75t_R register___U9742 ( .A(register__n11072), .Y(register__n6235) );
  BUFx2_ASAP7_75t_R register___U9743 ( .A(register__n6239), .Y(register__n6238) );
  BUFx2_ASAP7_75t_R register___U9744 ( .A(register__n12869), .Y(register__n6239) );
  BUFx2_ASAP7_75t_R register___U9745 ( .A(register__n6241), .Y(register__n6240) );
  BUFx2_ASAP7_75t_R register___U9746 ( .A(register__n13291), .Y(register__n6241) );
  BUFx2_ASAP7_75t_R register___U9747 ( .A(register__n6243), .Y(register__n6242) );
  BUFx2_ASAP7_75t_R register___U9748 ( .A(register__n12529), .Y(register__n6243) );
  BUFx2_ASAP7_75t_R register___U9749 ( .A(register__n6245), .Y(register__n6244) );
  BUFx2_ASAP7_75t_R register___U9750 ( .A(register__n12865), .Y(register__n6245) );
  BUFx2_ASAP7_75t_R register___U9751 ( .A(register__n13195), .Y(register__n6246) );
  BUFx2_ASAP7_75t_R register___U9752 ( .A(register__n13293), .Y(register__n6247) );
  BUFx2_ASAP7_75t_R register___U9753 ( .A(register__n6249), .Y(register__n6248) );
  BUFx2_ASAP7_75t_R register___U9754 ( .A(register__n6257), .Y(register__n6256) );
  BUFx2_ASAP7_75t_R register___U9755 ( .A(register__n13285), .Y(register__n6257) );
  BUFx2_ASAP7_75t_R register___U9756 ( .A(register__n6259), .Y(register__n6258) );
  OR2x2_ASAP7_75t_R register___U9757 ( .A(register__n6261), .B(register__n6262), .Y(register__n6260) );
  BUFx2_ASAP7_75t_R register___U9758 ( .A(register__n6987), .Y(register__n6261) );
  BUFx2_ASAP7_75t_R register___U9759 ( .A(register__n6988), .Y(register__n6262) );
  NOR2x1p5_ASAP7_75t_R register___U9760 ( .A(register__net89597), .B(register__n4920), .Y(register__n6987) );
  NOR2x1p5_ASAP7_75t_R register___U9761 ( .A(register__net64348), .B(register__n2220), .Y(register__n6988) );
  OR2x2_ASAP7_75t_R register___U9762 ( .A(register__n6264), .B(register__n8667), .Y(register__n6263) );
  BUFx2_ASAP7_75t_R register___U9763 ( .A(register__n8666), .Y(register__n6264) );
  NOR2x1p5_ASAP7_75t_R register___U9764 ( .A(register__net91219), .B(register__n1887), .Y(register__n8666) );
  BUFx12f_ASAP7_75t_R register___U9765 ( .A(register__n12450), .Y(register__n6268) );
  BUFx4f_ASAP7_75t_R register___U9766 ( .A(register__n6267), .Y(register__n12439) );
  BUFx4f_ASAP7_75t_R register___U9767 ( .A(register__net106240), .Y(register__net97246) );
  BUFx4f_ASAP7_75t_R register___U9768 ( .A(register__n7713), .Y(register__n8331) );
  BUFx3_ASAP7_75t_R register___U9769 ( .A(register__n6521), .Y(register__n6520) );
  BUFx3_ASAP7_75t_R register___U9770 ( .A(register__n6273), .Y(register__n6271) );
  BUFx4f_ASAP7_75t_R register___U9771 ( .A(register__n6273), .Y(register__n6272) );
  BUFx6f_ASAP7_75t_R register___U9772 ( .A(register__n6757), .Y(register__n6273) );
  BUFx4f_ASAP7_75t_R register___U9773 ( .A(register__n6271), .Y(register__n11181) );
  BUFx4f_ASAP7_75t_R register___U9774 ( .A(register__n6758), .Y(register__n6757) );
  BUFx3_ASAP7_75t_R register___U9775 ( .A(register__n6541), .Y(register__n6274) );
  BUFx3_ASAP7_75t_R register___U9776 ( .A(register__n7139), .Y(register__n6275) );
  BUFx3_ASAP7_75t_R register___U9777 ( .A(register__net103947), .Y(register__net114528) );
  BUFx4f_ASAP7_75t_R register___U9778 ( .A(register__net114528), .Y(register__net97186) );
  BUFx3_ASAP7_75t_R register___U9779 ( .A(register__n8108), .Y(register__n6276) );
  BUFx3_ASAP7_75t_R register___U9780 ( .A(register__n6525), .Y(register__n6277) );
  BUFx3_ASAP7_75t_R register___U9781 ( .A(register__n7388), .Y(register__n6278) );
  BUFx4f_ASAP7_75t_R register___U9782 ( .A(register__n6278), .Y(register__n8727) );
  BUFx3_ASAP7_75t_R register___U9783 ( .A(register__n6527), .Y(register__n6526) );
  BUFx3_ASAP7_75t_R register___U9784 ( .A(register__net112584), .Y(register__net114518) );
  BUFx3_ASAP7_75t_R register___U9785 ( .A(register__n6530), .Y(register__n6529) );
  BUFx3_ASAP7_75t_R register___U9786 ( .A(register__n8180), .Y(register__n6279) );
  BUFx3_ASAP7_75t_R register___U9787 ( .A(register__n6534), .Y(register__n6533) );
  BUFx3_ASAP7_75t_R register___U9788 ( .A(register__n8534), .Y(register__n6280) );
  BUFx3_ASAP7_75t_R register___U9789 ( .A(register__n7719), .Y(register__n6281) );
  BUFx3_ASAP7_75t_R register___U9790 ( .A(register__net90225), .Y(register__net114504) );
  BUFx2_ASAP7_75t_R register___U9791 ( .A(register__net90225), .Y(register__net114505) );
  BUFx12f_ASAP7_75t_R register___U9792 ( .A(register__n10336), .Y(register__n6282) );
  BUFx2_ASAP7_75t_R register___U9793 ( .A(Reg_data[470]), .Y(register__n6283) );
  BUFx3_ASAP7_75t_R register___U9794 ( .A(register__n10520), .Y(register__n6284) );
  BUFx2_ASAP7_75t_R register___U9795 ( .A(register__n10520), .Y(register__n6285) );
  BUFx4f_ASAP7_75t_R register___U9796 ( .A(register__n10520), .Y(register__n6286) );
  BUFx6f_ASAP7_75t_R register___U9797 ( .A(register__n10521), .Y(register__n10520) );
  BUFx4f_ASAP7_75t_R register___U9798 ( .A(register__n4956), .Y(register__n10521) );
  BUFx2_ASAP7_75t_R register___U9799 ( .A(Reg_data[400]), .Y(register__n6287) );
  BUFx6f_ASAP7_75t_R register___U9800 ( .A(register__n9410), .Y(register__n9409) );
  BUFx4f_ASAP7_75t_R register___U9801 ( .A(register__n5828), .Y(register__n9410) );
  BUFx2_ASAP7_75t_R register___U9802 ( .A(Reg_data[390]), .Y(register__net114451) );
  BUFx3_ASAP7_75t_R register___U9803 ( .A(register__net114452), .Y(register__net114453) );
  BUFx2_ASAP7_75t_R register___U9804 ( .A(Reg_data[384]), .Y(register__n6288) );
  BUFx6f_ASAP7_75t_R register___U9805 ( .A(register__n9412), .Y(register__n9411) );
  BUFx4f_ASAP7_75t_R register___U9806 ( .A(register__n5506), .Y(register__n9412) );
  BUFx3_ASAP7_75t_R register___U9807 ( .A(register__n6290), .Y(register__n6289) );
  BUFx2_ASAP7_75t_R register___U9808 ( .A(Reg_data[264]), .Y(register__n6290) );
  BUFx4f_ASAP7_75t_R register___U9809 ( .A(register__n6289), .Y(register__n8721) );
  BUFx3_ASAP7_75t_R register___U9810 ( .A(register__net114438), .Y(register__net114437) );
  BUFx2_ASAP7_75t_R register___U9811 ( .A(Reg_data[261]), .Y(register__net114438) );
  BUFx4f_ASAP7_75t_R register___U9812 ( .A(register__net114437), .Y(register__net97194) );
  BUFx3_ASAP7_75t_R register___U9813 ( .A(register__n6292), .Y(register__n6291) );
  BUFx2_ASAP7_75t_R register___U9814 ( .A(Reg_data[257]), .Y(register__n6292) );
  BUFx4f_ASAP7_75t_R register___U9815 ( .A(register__n6291), .Y(register__n7987) );
  BUFx2_ASAP7_75t_R register___U9816 ( .A(Reg_data[391]), .Y(register__n6293) );
  BUFx6f_ASAP7_75t_R register___U9817 ( .A(register__n9414), .Y(register__n9413) );
  BUFx4f_ASAP7_75t_R register___U9818 ( .A(register__n5653), .Y(register__n9414) );
  BUFx2_ASAP7_75t_R register___U9819 ( .A(Reg_data[252]), .Y(register__n6294) );
  BUFx6f_ASAP7_75t_R register___U9820 ( .A(register__n10154), .Y(register__n10153) );
  BUFx4f_ASAP7_75t_R register___U9821 ( .A(register__n5655), .Y(register__n10154) );
  BUFx2_ASAP7_75t_R register___U9822 ( .A(Reg_data[539]), .Y(register__n6295) );
  BUFx6f_ASAP7_75t_R register___U9823 ( .A(register__n8820), .Y(register__n8819) );
  BUFx4f_ASAP7_75t_R register___U9824 ( .A(register__n5656), .Y(register__n8820) );
  BUFx3_ASAP7_75t_R register___U9825 ( .A(register__n6297), .Y(register__n6296) );
  BUFx2_ASAP7_75t_R register___U9826 ( .A(Reg_data[265]), .Y(register__n6297) );
  BUFx4f_ASAP7_75t_R register___U9827 ( .A(register__n6296), .Y(register__n8737) );
  INVx1_ASAP7_75t_R register___U9828 ( .A(register__n10627), .Y(register__n6298) );
  INVx1_ASAP7_75t_R register___U9829 ( .A(register__n10691), .Y(register__n6299) );
  INVx1_ASAP7_75t_R register___U9830 ( .A(register__n10800), .Y(register__n6300) );
  BUFx3_ASAP7_75t_R register___U9831 ( .A(register__n6304), .Y(register__n6303) );
  BUFx2_ASAP7_75t_R register___U9832 ( .A(Reg_data[980]), .Y(register__n6304) );
  BUFx3_ASAP7_75t_R register___U9833 ( .A(register__net114311), .Y(register__net114310) );
  BUFx2_ASAP7_75t_R register___U9834 ( .A(Reg_data[761]), .Y(register__net114311) );
  BUFx3_ASAP7_75t_R register___U9835 ( .A(register__n6306), .Y(register__n6305) );
  BUFx2_ASAP7_75t_R register___U9836 ( .A(Reg_data[758]), .Y(register__n6306) );
  BUFx3_ASAP7_75t_R register___U9837 ( .A(register__n6308), .Y(register__n6307) );
  BUFx2_ASAP7_75t_R register___U9838 ( .A(Reg_data[738]), .Y(register__n6308) );
  BUFx3_ASAP7_75t_R register___U9839 ( .A(register__n6310), .Y(register__n6309) );
  BUFx2_ASAP7_75t_R register___U9840 ( .A(Reg_data[736]), .Y(register__n6310) );
  BUFx3_ASAP7_75t_R register___U9841 ( .A(register__n6312), .Y(register__n6311) );
  BUFx2_ASAP7_75t_R register___U9842 ( .A(Reg_data[720]), .Y(register__n6312) );
  BUFx3_ASAP7_75t_R register___U9843 ( .A(register__net114291), .Y(register__net114290) );
  BUFx2_ASAP7_75t_R register___U9844 ( .A(Reg_data[710]), .Y(register__net114291) );
  BUFx3_ASAP7_75t_R register___U9845 ( .A(register__n6314), .Y(register__n6313) );
  BUFx2_ASAP7_75t_R register___U9846 ( .A(Reg_data[707]), .Y(register__n6314) );
  BUFx3_ASAP7_75t_R register___U9847 ( .A(register__n6316), .Y(register__n6315) );
  BUFx2_ASAP7_75t_R register___U9848 ( .A(Reg_data[705]), .Y(register__n6316) );
  BUFx3_ASAP7_75t_R register___U9849 ( .A(register__n6318), .Y(register__n6317) );
  BUFx2_ASAP7_75t_R register___U9850 ( .A(Reg_data[692]), .Y(register__n6318) );
  BUFx3_ASAP7_75t_R register___U9851 ( .A(register__net114275), .Y(register__net114274) );
  BUFx2_ASAP7_75t_R register___U9852 ( .A(Reg_data[665]), .Y(register__net114275) );
  BUFx3_ASAP7_75t_R register___U9853 ( .A(register__n6320), .Y(register__n6319) );
  BUFx2_ASAP7_75t_R register___U9854 ( .A(Reg_data[642]), .Y(register__n6320) );
  BUFx3_ASAP7_75t_R register___U9855 ( .A(register__n9357), .Y(register__n6321) );
  BUFx2_ASAP7_75t_R register___U9856 ( .A(register__n9357), .Y(register__n6323) );
  BUFx3_ASAP7_75t_R register___U9857 ( .A(register__n6325), .Y(register__n6324) );
  BUFx2_ASAP7_75t_R register___U9858 ( .A(Reg_data[610]), .Y(register__n6325) );
  BUFx3_ASAP7_75t_R register___U9859 ( .A(register__n6327), .Y(register__n6326) );
  BUFx2_ASAP7_75t_R register___U9860 ( .A(Reg_data[530]), .Y(register__n6327) );
  BUFx3_ASAP7_75t_R register___U9861 ( .A(register__n6329), .Y(register__n6328) );
  BUFx2_ASAP7_75t_R register___U9862 ( .A(Reg_data[520]), .Y(register__n6329) );
  BUFx3_ASAP7_75t_R register___U9863 ( .A(register__net114249), .Y(register__net114248) );
  BUFx2_ASAP7_75t_R register___U9864 ( .A(Reg_data[517]), .Y(register__net114249) );
  BUFx3_ASAP7_75t_R register___U9865 ( .A(register__n6331), .Y(register__n6330) );
  BUFx2_ASAP7_75t_R register___U9866 ( .A(Reg_data[516]), .Y(register__n6331) );
  BUFx3_ASAP7_75t_R register___U9867 ( .A(register__n6333), .Y(register__n6332) );
  BUFx2_ASAP7_75t_R register___U9868 ( .A(Reg_data[513]), .Y(register__n6333) );
  BUFx3_ASAP7_75t_R register___U9869 ( .A(register__n6335), .Y(register__n6334) );
  BUFx2_ASAP7_75t_R register___U9870 ( .A(Reg_data[437]), .Y(register__n6335) );
  BUFx3_ASAP7_75t_R register___U9871 ( .A(register__n6337), .Y(register__n6336) );
  BUFx2_ASAP7_75t_R register___U9872 ( .A(Reg_data[424]), .Y(register__n6337) );
  BUFx3_ASAP7_75t_R register___U9873 ( .A(register__net114229), .Y(register__net114228) );
  BUFx2_ASAP7_75t_R register___U9874 ( .A(Reg_data[422]), .Y(register__net114229) );
  BUFx3_ASAP7_75t_R register___U9875 ( .A(register__net114225), .Y(register__net114224) );
  BUFx2_ASAP7_75t_R register___U9876 ( .A(Reg_data[421]), .Y(register__net114225) );
  BUFx3_ASAP7_75t_R register___U9877 ( .A(register__n6339), .Y(register__n6338) );
  BUFx2_ASAP7_75t_R register___U9878 ( .A(Reg_data[419]), .Y(register__n6339) );
  BUFx3_ASAP7_75t_R register___U9879 ( .A(register__n6341), .Y(register__n6340) );
  BUFx2_ASAP7_75t_R register___U9880 ( .A(Reg_data[387]), .Y(register__n6341) );
  BUFx3_ASAP7_75t_R register___U9881 ( .A(register__n6343), .Y(register__n6342) );
  BUFx2_ASAP7_75t_R register___U9882 ( .A(Reg_data[360]), .Y(register__n6343) );
  BUFx3_ASAP7_75t_R register___U9883 ( .A(register__net114209), .Y(register__net114208) );
  BUFx2_ASAP7_75t_R register___U9884 ( .A(Reg_data[971]), .Y(register__net114209) );
  BUFx3_ASAP7_75t_R register___U9885 ( .A(register__n6345), .Y(register__n6344) );
  BUFx2_ASAP7_75t_R register___U9886 ( .A(Reg_data[813]), .Y(register__n6345) );
  BUFx3_ASAP7_75t_R register___U9887 ( .A(register__net114201), .Y(register__net114200) );
  BUFx2_ASAP7_75t_R register___U9888 ( .A(Reg_data[970]), .Y(register__net114201) );
  BUFx3_ASAP7_75t_R register___U9889 ( .A(register__net114197), .Y(register__net114196) );
  BUFx2_ASAP7_75t_R register___U9890 ( .A(Reg_data[687]), .Y(register__net114197) );
  BUFx3_ASAP7_75t_R register___U9891 ( .A(register__n6347), .Y(register__n6346) );
  BUFx2_ASAP7_75t_R register___U9892 ( .A(Reg_data[638]), .Y(register__n6347) );
  BUFx3_ASAP7_75t_R register___U9893 ( .A(register__n6349), .Y(register__n6348) );
  BUFx2_ASAP7_75t_R register___U9894 ( .A(Reg_data[521]), .Y(register__n6349) );
  BUFx3_ASAP7_75t_R register___U9895 ( .A(register__n6351), .Y(register__n6350) );
  BUFx2_ASAP7_75t_R register___U9896 ( .A(Reg_data[423]), .Y(register__n6351) );
  BUFx3_ASAP7_75t_R register___U9897 ( .A(register__n6353), .Y(register__n6352) );
  BUFx2_ASAP7_75t_R register___U9898 ( .A(Reg_data[627]), .Y(register__n6353) );
  BUFx3_ASAP7_75t_R register___U9899 ( .A(register__n6355), .Y(register__n6354) );
  BUFx2_ASAP7_75t_R register___U9900 ( .A(Reg_data[823]), .Y(register__n6355) );
  BUFx3_ASAP7_75t_R register___U9901 ( .A(register__n6357), .Y(register__n6356) );
  BUFx2_ASAP7_75t_R register___U9902 ( .A(Reg_data[46]), .Y(register__n6357) );
  BUFx3_ASAP7_75t_R register___U9903 ( .A(register__net114169), .Y(register__net114168) );
  BUFx2_ASAP7_75t_R register___U9904 ( .A(Reg_data[810]), .Y(register__net114169) );
  BUFx3_ASAP7_75t_R register___U9905 ( .A(register__n6359), .Y(register__n6358) );
  BUFx2_ASAP7_75t_R register___U9906 ( .A(Reg_data[979]), .Y(register__n6359) );
  BUFx3_ASAP7_75t_R register___U9907 ( .A(register__n6361), .Y(register__n6360) );
  BUFx2_ASAP7_75t_R register___U9908 ( .A(Reg_data[983]), .Y(register__n6361) );
  BUFx3_ASAP7_75t_R register___U9909 ( .A(register__n6363), .Y(register__n6362) );
  BUFx2_ASAP7_75t_R register___U9910 ( .A(Reg_data[972]), .Y(register__n6363) );
  BUFx3_ASAP7_75t_R register___U9911 ( .A(register__n6365), .Y(register__n6364) );
  BUFx2_ASAP7_75t_R register___U9912 ( .A(Reg_data[205]), .Y(register__n6365) );
  BUFx12f_ASAP7_75t_R register___U9913 ( .A(register__n10125), .Y(register__n6366) );
  BUFx12f_ASAP7_75t_R register___U9914 ( .A(register__n6366), .Y(register__n10124) );
  BUFx3_ASAP7_75t_R register___U9915 ( .A(register__n6368), .Y(register__n6367) );
  BUFx2_ASAP7_75t_R register___U9916 ( .A(Reg_data[236]), .Y(register__n6368) );
  BUFx3_ASAP7_75t_R register___U9917 ( .A(register__n6370), .Y(register__n6369) );
  BUFx2_ASAP7_75t_R register___U9918 ( .A(Reg_data[439]), .Y(register__n6370) );
  BUFx3_ASAP7_75t_R register___U9919 ( .A(register__n6372), .Y(register__n6371) );
  BUFx2_ASAP7_75t_R register___U9920 ( .A(Reg_data[489]), .Y(register__n6372) );
  BUFx3_ASAP7_75t_R register___U9921 ( .A(register__n6374), .Y(register__n6373) );
  BUFx2_ASAP7_75t_R register___U9922 ( .A(Reg_data[543]), .Y(register__n6374) );
  BUFx2_ASAP7_75t_R register___U9923 ( .A(register__n10171), .Y(register__n6375) );
  BUFx2_ASAP7_75t_R register___U9924 ( .A(register__n10171), .Y(register__n6376) );
  BUFx4f_ASAP7_75t_R register___U9925 ( .A(register__n10171), .Y(register__n6377) );
  BUFx3_ASAP7_75t_R register___U9926 ( .A(register__n6379), .Y(register__n6378) );
  BUFx2_ASAP7_75t_R register___U9927 ( .A(Reg_data[575]), .Y(register__n6379) );
  BUFx3_ASAP7_75t_R register___U9928 ( .A(register__net114120), .Y(register__net114119) );
  BUFx2_ASAP7_75t_R register___U9929 ( .A(Reg_data[504]), .Y(register__net114120) );
  BUFx3_ASAP7_75t_R register___U9930 ( .A(register__net114110), .Y(register__net114109) );
  BUFx2_ASAP7_75t_R register___U9931 ( .A(Reg_data[399]), .Y(register__net114110) );
  BUFx2_ASAP7_75t_R register___U9932 ( .A(register__net90525), .Y(register__net114112) );
  BUFx4f_ASAP7_75t_R register___U9933 ( .A(register__net90525), .Y(register__net114113) );
  BUFx3_ASAP7_75t_R register___U9934 ( .A(register__n6381), .Y(register__n6380) );
  BUFx2_ASAP7_75t_R register___U9935 ( .A(Reg_data[766]), .Y(register__n6381) );
  BUFx3_ASAP7_75t_R register___U9936 ( .A(register__n6383), .Y(register__n6382) );
  BUFx2_ASAP7_75t_R register___U9937 ( .A(Reg_data[526]), .Y(register__n6383) );
  BUFx2_ASAP7_75t_R register___U9938 ( .A(register__n10208), .Y(register__n6384) );
  BUFx6f_ASAP7_75t_R register___U9939 ( .A(register__n10208), .Y(register__n6385) );
  BUFx3_ASAP7_75t_R register___U9940 ( .A(register__net114094), .Y(register__net114093) );
  BUFx2_ASAP7_75t_R register___U9941 ( .A(Reg_data[426]), .Y(register__net114094) );
  BUFx3_ASAP7_75t_R register___U9942 ( .A(register__n6387), .Y(register__n6386) );
  BUFx2_ASAP7_75t_R register___U9943 ( .A(Reg_data[635]), .Y(register__n6387) );
  BUFx3_ASAP7_75t_R register___U9944 ( .A(register__n6389), .Y(register__n6388) );
  BUFx2_ASAP7_75t_R register___U9945 ( .A(Reg_data[689]), .Y(register__n6389) );
  BUFx3_ASAP7_75t_R register___U9946 ( .A(register__n6391), .Y(register__n6390) );
  BUFx2_ASAP7_75t_R register___U9947 ( .A(Reg_data[251]), .Y(register__n6391) );
  BUFx3_ASAP7_75t_R register___U9948 ( .A(register__n6393), .Y(register__n6392) );
  BUFx2_ASAP7_75t_R register___U9949 ( .A(Reg_data[319]), .Y(register__n6393) );
  BUFx12f_ASAP7_75t_R register___U9950 ( .A(register__n3377), .Y(register__n12133) );
  BUFx12f_ASAP7_75t_R register___U9951 ( .A(register__n6680), .Y(register__n12138) );
  OA22x2_ASAP7_75t_R register___U9952 ( .A1(register__n12151), .A2(register__n2220), .B1(register__n10152), .B2(register__n3414), 
        .Y(register__n12789) );
  INVx1_ASAP7_75t_R register___U9953 ( .A(register__n3901), .Y(register__n6396) );
  OA22x2_ASAP7_75t_R register___U9954 ( .A1(register__n12226), .A2(register__n399), .B1(register__n10175), .B2(register__n3380), 
        .Y(register__n13299) );
  OA22x2_ASAP7_75t_R register___U9955 ( .A1(register__net64356), .A2(register__n7327), .B1(register__net90717), .B2(
        n11831), .Y(register__n12568) );
  OA22x2_ASAP7_75t_R register___U9956 ( .A1(register__net64670), .A2(register__n996), .B1(register__n10164), .B2(register__n969), 
        .Y(register__n13201) );
  INVx1_ASAP7_75t_R register___U9957 ( .A(register__n4080), .Y(register__n6399) );
  OA22x2_ASAP7_75t_R register___U9958 ( .A1(register__n12280), .A2(register__n399), .B1(register__n10235), .B2(register__n3606), 
        .Y(register__n13297) );
  INVx1_ASAP7_75t_R register___U9959 ( .A(register__n4886), .Y(register__n6400) );
  OA22x2_ASAP7_75t_R register___U9960 ( .A1(register__net63326), .A2(register__n977), .B1(register__n10271), .B2(register__n974), 
        .Y(register__n13185) );
  OA22x2_ASAP7_75t_R register___U9961 ( .A1(register__n12313), .A2(register__n988), .B1(register__n7488), .B2(register__n971), 
        .Y(register__n13188) );
  INVx1_ASAP7_75t_R register___U9962 ( .A(register__n5781), .Y(register__n6401) );
  OA22x2_ASAP7_75t_R register___U9963 ( .A1(register__net64418), .A2(register__n1004), .B1(register__net107944), .B2(
        n973), .Y(register__n13198) );
  INVx1_ASAP7_75t_R register___U9964 ( .A(register__n5787), .Y(register__n6402) );
  OA22x2_ASAP7_75t_R register___U9965 ( .A1(register__net64420), .A2(register__n103), .B1(register__net103925), .B2(
        n1146), .Y(register__n13166) );
  INVx2_ASAP7_75t_R register___U9966 ( .A(register__n12471), .Y(register__n12456) );
  BUFx4f_ASAP7_75t_R register___U9967 ( .A(register__n3214), .Y(register__n12471) );
  INVx2_ASAP7_75t_R register___U9968 ( .A(register__n9406), .Y(register__n11964) );
  BUFx6f_ASAP7_75t_R register___U9969 ( .A(register__n4650), .Y(register__n12213) );
  BUFx6f_ASAP7_75t_R register___U9970 ( .A(register__n4649), .Y(register__n12211) );
  BUFx6f_ASAP7_75t_R register___U9971 ( .A(register__n6405), .Y(register__n12013) );
  BUFx6f_ASAP7_75t_R register___U9972 ( .A(register__n6405), .Y(register__n12014) );
  BUFx6f_ASAP7_75t_R register___U9973 ( .A(register__n6405), .Y(register__n12007) );
  BUFx4f_ASAP7_75t_R register___U9974 ( .A(register__n6405), .Y(register__n12010) );
  BUFx4f_ASAP7_75t_R register___U9975 ( .A(register__n6405), .Y(register__n12009) );
  BUFx6f_ASAP7_75t_R register___U9976 ( .A(register__net139023), .Y(register__net63038) );
  BUFx6f_ASAP7_75t_R register___U9977 ( .A(register__net129690), .Y(register__net63032) );
  INVx1_ASAP7_75t_R register___U9978 ( .A(register__n4019), .Y(register__n6408) );
  INVx1_ASAP7_75t_R register___U9979 ( .A(register__n4450), .Y(register__n6409) );
  INVx1_ASAP7_75t_R register___U9980 ( .A(register__n4452), .Y(register__n6410) );
  INVx1_ASAP7_75t_R register___U9981 ( .A(register__n4454), .Y(register__n6411) );
  AND4x1_ASAP7_75t_R register___U9982 ( .A(register__n6411), .B(register__n6409), .C(register__n8560), .D(register__n4453), .Y(
        n10950) );
  INVx1_ASAP7_75t_R register___U9983 ( .A(register__n3880), .Y(register__n6412) );
  INVx1_ASAP7_75t_R register___U9984 ( .A(register__n4310), .Y(register__n6413) );
  INVx1_ASAP7_75t_R register___U9985 ( .A(register__n4312), .Y(register__n6414) );
  INVx1_ASAP7_75t_R register___U9986 ( .A(register__n4315), .Y(register__n6415) );
  INVx1_ASAP7_75t_R register___U9987 ( .A(register__n5582), .Y(register__n6416) );
  INVx1_ASAP7_75t_R register___U9988 ( .A(register__n5279), .Y(register__n6417) );
  INVx1_ASAP7_75t_R register___U9989 ( .A(register__n5282), .Y(register__n6418) );
  AND4x1_ASAP7_75t_R register___U9990 ( .A(register__n1298), .B(register__n8256), .C(register__n6418), .D(register__n5281), .Y(
        n10611) );
  INVx1_ASAP7_75t_R register___U9991 ( .A(register__n4353), .Y(register__n6421) );
  INVx1_ASAP7_75t_R register___U9992 ( .A(register__n4356), .Y(register__n6422) );
  INVx1_ASAP7_75t_R register___U9993 ( .A(register__n4357), .Y(register__n6423) );
  INVx1_ASAP7_75t_R register___U9994 ( .A(register__n11092), .Y(register__n6427) );
  INVx1_ASAP7_75t_R register___U9995 ( .A(register__n4713), .Y(register__n6428) );
  INVx1_ASAP7_75t_R register___U9996 ( .A(register__n4715), .Y(register__n6429) );
  OA22x2_ASAP7_75t_R register___U9997 ( .A1(register__net63996), .A2(register__n1137), .B1(register__net103941), .B2(
        n1143), .Y(register__n13162) );
  OA22x2_ASAP7_75t_R register___U9998 ( .A1(register__n11935), .A2(register__n4033), .B1(register__n9577), .B2(register__n3329), 
        .Y(register__n12552) );
  OA22x2_ASAP7_75t_R register___U9999 ( .A1(register__n12031), .A2(register__n7327), .B1(register__n5174), .B2(register__n5525), 
        .Y(register__n12575) );
  INVx1_ASAP7_75t_R register___U10000 ( .A(register__n4391), .Y(register__n6432) );
  OA22x2_ASAP7_75t_R register___U10001 ( .A1(register__net63164), .A2(register__n955), .B1(register__net90925), .B2(
        n960), .Y(register__n13015) );
  OA22x2_ASAP7_75t_R register___U10002 ( .A1(register__n12314), .A2(register__n1137), .B1(register__n9211), .B2(register__n1148), 
        .Y(register__n13158) );
  OA22x2_ASAP7_75t_R register___U10003 ( .A1(register__net64924), .A2(register__n103), .B1(register__n8722), .B2(register__n1145), 
        .Y(register__n13172) );
  OA22x2_ASAP7_75t_R register___U10004 ( .A1(register__net64352), .A2(register__n3022), .B1(register__net91375), .B2(
        n1585), .Y(register__n12707) );
  OA22x2_ASAP7_75t_R register___U10005 ( .A1(register__n12153), .A2(register__n3022), .B1(register__n9505), .B2(register__n1584), 
        .Y(register__n12705) );
  OA22x2_ASAP7_75t_R register___U10006 ( .A1(register__n12152), .A2(register__n2803), .B1(register__n2982), .B2(register__n9509), 
        .Y(register__n12875) );
  OA22x2_ASAP7_75t_R register___U10007 ( .A1(register__net62678), .A2(register__n4033), .B1(register__n8797), .B2(
        n11843), .Y(register__n12522) );
  INVx1_ASAP7_75t_R register___U10008 ( .A(register__n5771), .Y(register__n6438) );
  OA22x2_ASAP7_75t_R register___U10009 ( .A1(register__n3443), .A2(register__n103), .B1(register__n7661), .B2(register__n1058), 
        .Y(register__n13161) );
  INVx1_ASAP7_75t_R register___U10010 ( .A(register__n3960), .Y(register__n6439) );
  OA22x2_ASAP7_75t_R register___U10011 ( .A1(register__net62824), .A2(register__n1140), .B1(register__net91255), .B2(
        n1146), .Y(register__n13150) );
  OA22x2_ASAP7_75t_R register___U10012 ( .A1(register__net64004), .A2(register__n951), .B1(register__net90521), .B2(
        n960), .Y(register__n13024) );
  OA22x2_ASAP7_75t_R register___U10013 ( .A1(register__n12397), .A2(register__n1139), .B1(register__n9565), .B2(register__n1143), 
        .Y(register__n13153) );
  OA22x2_ASAP7_75t_R register___U10014 ( .A1(register__n12281), .A2(register__n1049), .B1(register__n10241), .B2(register__n3908), 
        .Y(register__n13272) );
  OA22x2_ASAP7_75t_R register___U10015 ( .A1(register__n12292), .A2(register__n105), .B1(register__n7999), .B2(register__n1669), 
        .Y(register__n12644) );
  INVx1_ASAP7_75t_R register___U10016 ( .A(register__n3744), .Y(register__n6442) );
  BUFx12f_ASAP7_75t_R register___U10017 ( .A(register__net73061), .Y(register__net73059) );
  OA22x2_ASAP7_75t_R register___U10018 ( .A1(register__net63328), .A2(register__n1137), .B1(register__n9213), .B2(register__n1145), .Y(register__n13155) );
  OA22x2_ASAP7_75t_R register___U10019 ( .A1(register__n12231), .A2(register__n1917), .B1(register__n10311), .B2(register__n2135), 
        .Y(register__n12902) );
  OA22x2_ASAP7_75t_R register___U10020 ( .A1(register__n99), .A2(register__n576), .B1(register__n10319), .B2(register__n580), .Y(
        n13221) );
  INVx1_ASAP7_75t_R register___U10021 ( .A(register__n4537), .Y(register__n6444) );
  OA22x2_ASAP7_75t_R register___U10022 ( .A1(register__n12197), .A2(register__n952), .B1(register__n9333), .B2(register__n959), 
        .Y(register__n13023) );
  OA22x2_ASAP7_75t_R register___U10023 ( .A1(register__net64776), .A2(register__n7327), .B1(register__net116359), .B2(
        n5172), .Y(register__n12572) );
  INVx1_ASAP7_75t_R register___U10024 ( .A(register__n4597), .Y(register__n6446) );
  INVx1_ASAP7_75t_R register___U10025 ( .A(register__n11004), .Y(register__n6447) );
  INVx1_ASAP7_75t_R register___U10026 ( .A(register__n3000), .Y(register__n6449) );
  INVx1_ASAP7_75t_R register___U10027 ( .A(register__n3132), .Y(register__n6450) );
  INVx1_ASAP7_75t_R register___U10028 ( .A(register__n3135), .Y(register__n6452) );
  INVx1_ASAP7_75t_R register___U10029 ( .A(register__n3619), .Y(register__n6454) );
  INVx1_ASAP7_75t_R register___U10030 ( .A(register__n3621), .Y(register__n6455) );
  INVx1_ASAP7_75t_R register___U10031 ( .A(register__n3622), .Y(register__n6456) );
  INVx1_ASAP7_75t_R register___U10032 ( .A(register__n3624), .Y(register__n6458) );
  INVx1_ASAP7_75t_R register___U10033 ( .A(register__n3626), .Y(register__n6459) );
  OA22x2_ASAP7_75t_R register___U10034 ( .A1(register__n12347), .A2(register__n11816), .B1(register__n9445), .B2(register__n1592), 
        .Y(register__n12699) );
  OA22x2_ASAP7_75t_R register___U10035 ( .A1(register__n12255), .A2(register__n1137), .B1(register__n9479), .B2(register__n1148), 
        .Y(register__n13160) );
  INVx1_ASAP7_75t_R register___U10036 ( .A(register__n3740), .Y(register__n6460) );
  INVx2_ASAP7_75t_R register___U10037 ( .A(register__n12037), .Y(register__n12022) );
  OA22x2_ASAP7_75t_R register___U10038 ( .A1(register__n3442), .A2(register__n1139), .B1(register__n9485), .B2(register__n1141), 
        .Y(register__n13176) );
  OA22x2_ASAP7_75t_R register___U10039 ( .A1(register__net63244), .A2(register__n1755), .B1(register__net90637), .B2(
        n3821), .Y(register__n13123) );
  INVx1_ASAP7_75t_R register___U10040 ( .A(register__n2989), .Y(register__n6461) );
  OA22x2_ASAP7_75t_R register___U10041 ( .A1(register__net64664), .A2(register__n3719), .B1(register__n10379), .B2(
        n1163), .Y(register__n13382) );
  BUFx12f_ASAP7_75t_R register___U10042 ( .A(register__n3308), .Y(register__n6462) );
  BUFx12f_ASAP7_75t_R register___U10043 ( .A(register__n11815), .Y(register__n11814) );
  BUFx2_ASAP7_75t_R register___U10044 ( .A(register__n10664), .Y(register__n6470) );
  INVx2_ASAP7_75t_R register___U10045 ( .A(register__n10343), .Y(register__n11227) );
  INVx2_ASAP7_75t_R register___U10046 ( .A(register__net93375), .Y(register__C6423_net61304) );
  BUFx2_ASAP7_75t_R register___U10047 ( .A(register__n10893), .Y(register__n6471) );
  BUFx2_ASAP7_75t_R register___U10048 ( .A(register__n11415), .Y(register__n6472) );
  INVx2_ASAP7_75t_R register___U10049 ( .A(register__net88813), .Y(register__C6423_net61194) );
  BUFx2_ASAP7_75t_R register___U10050 ( .A(register__n11547), .Y(register__n6474) );
  BUFx2_ASAP7_75t_R register___U10051 ( .A(register__n11106), .Y(register__n6475) );
  BUFx2_ASAP7_75t_R register___U10052 ( .A(register__n11351), .Y(register__n6476) );
  BUFx2_ASAP7_75t_R register___U10053 ( .A(register__n11457), .Y(register__n6477) );
  INVx2_ASAP7_75t_R register___U10054 ( .A(register__n10393), .Y(register__n11063) );
  BUFx2_ASAP7_75t_R register___U10055 ( .A(register__n10788), .Y(register__n6478) );
  BUFx2_ASAP7_75t_R register___U10056 ( .A(register__n11502), .Y(register__n6479) );
  INVx2_ASAP7_75t_R register___U10057 ( .A(register__n10413), .Y(register__n11043) );
  BUFx2_ASAP7_75t_R register___U10058 ( .A(register__n10934), .Y(register__n6480) );
  BUFx2_ASAP7_75t_R register___U10059 ( .A(register__n10869), .Y(register__n6481) );
  BUFx2_ASAP7_75t_R register___U10060 ( .A(register__n11304), .Y(register__n6482) );
  INVx2_ASAP7_75t_R register___U10061 ( .A(register__n9475), .Y(register__n10957) );
  INVx2_ASAP7_75t_R register___U10062 ( .A(register__n9449), .Y(register__n10867) );
  BUFx2_ASAP7_75t_R register___U10063 ( .A(register__n11434), .Y(register__n6483) );
  BUFx2_ASAP7_75t_R register___U10064 ( .A(register__n11180), .Y(register__n6484) );
  INVx2_ASAP7_75t_R register___U10065 ( .A(register__n9465), .Y(register__n11435) );
  BUFx2_ASAP7_75t_R register___U10066 ( .A(register__C6422_net60219), .Y(register__net113240) );
  BUFx2_ASAP7_75t_R register___U10067 ( .A(register__n10913), .Y(register__n6485) );
  BUFx2_ASAP7_75t_R register___U10068 ( .A(register__n10574), .Y(register__n6486) );
  BUFx2_ASAP7_75t_R register___U10069 ( .A(register__n10955), .Y(register__n6487) );
  BUFx2_ASAP7_75t_R register___U10070 ( .A(register__n10554), .Y(register__n6488) );
  BUFx2_ASAP7_75t_R register___U10071 ( .A(register__C6422_net59829), .Y(register__net113227) );
  INVx2_ASAP7_75t_R register___U10072 ( .A(register__n9543), .Y(register__n11454) );
  INVx2_ASAP7_75t_R register___U10073 ( .A(register__n9569), .Y(register__n11350) );
  INVx2_ASAP7_75t_R register___U10074 ( .A(register__n9511), .Y(register__n11305) );
  INVx2_ASAP7_75t_R register___U10075 ( .A(register__n9567), .Y(register__n11372) );
  BUFx2_ASAP7_75t_R register___U10076 ( .A(register__n11625), .Y(register__n6489) );
  BUFx2_ASAP7_75t_R register___U10077 ( .A(register__n11017), .Y(register__n6490) );
  BUFx2_ASAP7_75t_R register___U10078 ( .A(register__n11685), .Y(register__n6491) );
  BUFx2_ASAP7_75t_R register___U10079 ( .A(register__n11371), .Y(register__n6492) );
  BUFx2_ASAP7_75t_R register___U10080 ( .A(register__net94613), .Y(register__net113158) );
  BUFx4f_ASAP7_75t_R register___U10081 ( .A(register__net94613), .Y(register__net113159) );
  BUFx2_ASAP7_75t_R register___U10082 ( .A(register__net94610), .Y(register__net113150) );
  BUFx2_ASAP7_75t_R register___U10083 ( .A(register__n6501), .Y(register__n6500) );
  BUFx2_ASAP7_75t_R register___U10084 ( .A(register__n13303), .Y(register__n6501) );
  BUFx2_ASAP7_75t_R register___U10085 ( .A(register__n6503), .Y(register__n6502) );
  BUFx2_ASAP7_75t_R register___U10086 ( .A(register__n12543), .Y(register__n6503) );
  BUFx2_ASAP7_75t_R register___U10087 ( .A(register__n6505), .Y(register__n6504) );
  BUFx2_ASAP7_75t_R register___U10088 ( .A(register__n12545), .Y(register__n6505) );
  BUFx2_ASAP7_75t_R register___U10089 ( .A(register__n6511), .Y(register__n6510) );
  BUFx2_ASAP7_75t_R register___U10090 ( .A(register__n13287), .Y(register__n6511) );
  BUFx2_ASAP7_75t_R register___U10091 ( .A(register__n6513), .Y(register__n6512) );
  BUFx2_ASAP7_75t_R register___U10092 ( .A(register__n12822), .Y(register__n6513) );
  BUFx2_ASAP7_75t_R register___U10093 ( .A(register__n9390), .Y(register__n6514) );
  BUFx2_ASAP7_75t_R register___U10094 ( .A(register__n12533), .Y(register__n6515) );
  BUFx3_ASAP7_75t_R register___U10095 ( .A(register__n6517), .Y(register__n6516) );
  BUFx2_ASAP7_75t_R register___U10096 ( .A(register__n10903), .Y(register__n6517) );
  BUFx3_ASAP7_75t_R register___U10097 ( .A(register__n6519), .Y(register__n6518) );
  BUFx2_ASAP7_75t_R register___U10098 ( .A(register__n10904), .Y(register__n6519) );
  BUFx12f_ASAP7_75t_R register___U10099 ( .A(register__net99590), .Y(register__net112763) );
  BUFx12f_ASAP7_75t_R register___U10100 ( .A(register__net116957), .Y(register__net112764) );
  BUFx3_ASAP7_75t_R register___U10101 ( .A(register__n6807), .Y(register__n6806) );
  BUFx3_ASAP7_75t_R register___U10102 ( .A(register__net110255), .Y(register__net112748) );
  BUFx2_ASAP7_75t_R register___U10103 ( .A(Reg_data[784]), .Y(register__n6521) );
  BUFx6f_ASAP7_75t_R register___U10104 ( .A(register__n7329), .Y(register__n7328) );
  BUFx4f_ASAP7_75t_R register___U10105 ( .A(register__n6520), .Y(register__n7329) );
  BUFx3_ASAP7_75t_R register___U10106 ( .A(register__n8027), .Y(register__n6522) );
  BUFx4f_ASAP7_75t_R register___U10107 ( .A(register__n6522), .Y(register__n8711) );
  BUFx3_ASAP7_75t_R register___U10108 ( .A(register__net101470), .Y(register__net112736) );
  BUFx4f_ASAP7_75t_R register___U10109 ( .A(register__net112736), .Y(register__net97226) );
  BUFx12f_ASAP7_75t_R register___U10110 ( .A(register__n9675), .Y(register__n6523) );
  BUFx4f_ASAP7_75t_R register___U10111 ( .A(register__net89913), .Y(register__net112729) );
  BUFx2_ASAP7_75t_R register___U10112 ( .A(register__net89913), .Y(register__net112730) );
  BUFx3_ASAP7_75t_R register___U10113 ( .A(register__n8090), .Y(register__n6524) );
  BUFx12f_ASAP7_75t_R register___U10114 ( .A(register__net89598), .Y(register__net112724) );
  BUFx2_ASAP7_75t_R register___U10115 ( .A(Reg_data[583]), .Y(register__n6525) );
  BUFx6f_ASAP7_75t_R register___U10116 ( .A(register__n8689), .Y(register__n8688) );
  BUFx4f_ASAP7_75t_R register___U10117 ( .A(register__n6277), .Y(register__n8689) );
  BUFx2_ASAP7_75t_R register___U10118 ( .A(Reg_data[777]), .Y(register__n6527) );
  BUFx6f_ASAP7_75t_R register___U10119 ( .A(register__n7331), .Y(register__n7330) );
  BUFx4f_ASAP7_75t_R register___U10120 ( .A(register__n6526), .Y(register__n7331) );
  BUFx3_ASAP7_75t_R register___U10121 ( .A(register__n7195), .Y(register__n6528) );
  BUFx2_ASAP7_75t_R register___U10122 ( .A(Reg_data[780]), .Y(register__n6530) );
  BUFx6f_ASAP7_75t_R register___U10123 ( .A(register__n7333), .Y(register__n7332) );
  BUFx4f_ASAP7_75t_R register___U10124 ( .A(register__n6529), .Y(register__n7333) );
  BUFx3_ASAP7_75t_R register___U10125 ( .A(register__n7716), .Y(register__n6531) );
  BUFx3_ASAP7_75t_R register___U10126 ( .A(register__n9101), .Y(register__n6532) );
  BUFx2_ASAP7_75t_R register___U10127 ( .A(Reg_data[794]), .Y(register__n6534) );
  BUFx6f_ASAP7_75t_R register___U10128 ( .A(register__n7335), .Y(register__n7334) );
  BUFx4f_ASAP7_75t_R register___U10129 ( .A(register__n6533), .Y(register__n7335) );
  BUFx3_ASAP7_75t_R register___U10130 ( .A(register__n8190), .Y(register__n6535) );
  BUFx3_ASAP7_75t_R register___U10131 ( .A(register__net112639), .Y(register__net112638) );
  BUFx2_ASAP7_75t_R register___U10132 ( .A(Reg_data[601]), .Y(register__net112639) );
  BUFx4f_ASAP7_75t_R register___U10133 ( .A(register__net112638), .Y(register__net97238) );
  BUFx3_ASAP7_75t_R register___U10134 ( .A(register__n6537), .Y(register__n6536) );
  BUFx2_ASAP7_75t_R register___U10135 ( .A(Reg_data[594]), .Y(register__n6537) );
  BUFx4f_ASAP7_75t_R register___U10136 ( .A(register__n6536), .Y(register__n8709) );
  BUFx3_ASAP7_75t_R register___U10137 ( .A(register__n6539), .Y(register__n6538) );
  BUFx2_ASAP7_75t_R register___U10138 ( .A(Reg_data[580]), .Y(register__n6539) );
  BUFx4f_ASAP7_75t_R register___U10139 ( .A(register__n6538), .Y(register__n8713) );
  BUFx2_ASAP7_75t_R register___U10140 ( .A(Reg_data[432]), .Y(register__n6540) );
  BUFx6f_ASAP7_75t_R register___U10141 ( .A(register__n9334), .Y(register__n9333) );
  BUFx4f_ASAP7_75t_R register___U10142 ( .A(register__n6037), .Y(register__n9334) );
  BUFx2_ASAP7_75t_R register___U10143 ( .A(Reg_data[53]), .Y(register__n6541) );
  BUFx6f_ASAP7_75t_R register___U10144 ( .A(register__n10075), .Y(register__n10074) );
  BUFx4f_ASAP7_75t_R register___U10145 ( .A(register__n6274), .Y(register__n10075) );
  BUFx3_ASAP7_75t_R register___U10146 ( .A(register__net112616), .Y(register__net112615) );
  BUFx2_ASAP7_75t_R register___U10147 ( .A(Reg_data[331]), .Y(register__net112616) );
  BUFx4f_ASAP7_75t_R register___U10148 ( .A(register__net112615), .Y(register__net97182) );
  BUFx3_ASAP7_75t_R register___U10149 ( .A(register__n6543), .Y(register__n6542) );
  BUFx2_ASAP7_75t_R register___U10150 ( .A(Reg_data[599]), .Y(register__n6543) );
  BUFx4f_ASAP7_75t_R register___U10151 ( .A(register__n6542), .Y(register__n8725) );
  BUFx2_ASAP7_75t_R register___U10152 ( .A(Reg_data[540]), .Y(register__n6544) );
  BUFx6f_ASAP7_75t_R register___U10153 ( .A(register__n10137), .Y(register__n10136) );
  BUFx4f_ASAP7_75t_R register___U10154 ( .A(register__n5654), .Y(register__n10137) );
  BUFx2_ASAP7_75t_R register___U10155 ( .A(Reg_data[250]), .Y(register__n6545) );
  BUFx6f_ASAP7_75t_R register___U10156 ( .A(register__n10166), .Y(register__n10165) );
  BUFx4f_ASAP7_75t_R register___U10157 ( .A(register__n6042), .Y(register__n10166) );
  BUFx2_ASAP7_75t_R register___U10158 ( .A(Reg_data[253]), .Y(register__net112592) );
  BUFx2_ASAP7_75t_R register___U10159 ( .A(register__net89441), .Y(register__net112594) );
  BUFx4f_ASAP7_75t_R register___U10160 ( .A(register__net118023), .Y(register__net89441) );
  BUFx2_ASAP7_75t_R register___U10161 ( .A(Reg_data[591]), .Y(register__net112584) );
  BUFx6f_ASAP7_75t_R register___U10162 ( .A(register__net97157), .Y(register__net112585) );
  BUFx6f_ASAP7_75t_R register___U10163 ( .A(register__net97158), .Y(register__net97157) );
  BUFx4f_ASAP7_75t_R register___U10164 ( .A(register__net114518), .Y(register__net97158) );
  BUFx12f_ASAP7_75t_R register___U10165 ( .A(register__net112580), .Y(register__net112578) );
  INVx1_ASAP7_75t_R register___U10166 ( .A(register__n5553), .Y(register__n6546) );
  INVx1_ASAP7_75t_R register___U10167 ( .A(register__n11464), .Y(register__n6548) );
  INVx1_ASAP7_75t_R register___U10168 ( .A(register__n5599), .Y(register__n6549) );
  BUFx3_ASAP7_75t_R register___U10169 ( .A(register__net112550), .Y(register__net112549) );
  BUFx2_ASAP7_75t_R register___U10170 ( .A(Reg_data[805]), .Y(register__net112550) );
  BUFx3_ASAP7_75t_R register___U10171 ( .A(register__n6551), .Y(register__n6550) );
  BUFx2_ASAP7_75t_R register___U10172 ( .A(Reg_data[804]), .Y(register__n6551) );
  BUFx3_ASAP7_75t_R register___U10173 ( .A(register__net112542), .Y(register__net112541) );
  BUFx2_ASAP7_75t_R register___U10174 ( .A(Reg_data[741]), .Y(register__net112542) );
  BUFx3_ASAP7_75t_R register___U10175 ( .A(register__n6553), .Y(register__n6552) );
  BUFx2_ASAP7_75t_R register___U10176 ( .A(Reg_data[740]), .Y(register__n6553) );
  BUFx3_ASAP7_75t_R register___U10177 ( .A(register__net112534), .Y(register__net112533) );
  BUFx2_ASAP7_75t_R register___U10178 ( .A(Reg_data[697]), .Y(register__net112534) );
  BUFx3_ASAP7_75t_R register___U10179 ( .A(register__n6555), .Y(register__n6554) );
  BUFx2_ASAP7_75t_R register___U10180 ( .A(Reg_data[694]), .Y(register__n6555) );
  BUFx3_ASAP7_75t_R register___U10181 ( .A(register__n6557), .Y(register__n6556) );
  BUFx2_ASAP7_75t_R register___U10182 ( .A(Reg_data[672]), .Y(register__n6557) );
  BUFx3_ASAP7_75t_R register___U10183 ( .A(register__n6559), .Y(register__n6558) );
  BUFx2_ASAP7_75t_R register___U10184 ( .A(Reg_data[662]), .Y(register__n6559) );
  BUFx3_ASAP7_75t_R register___U10185 ( .A(register__n6561), .Y(register__n6560) );
  BUFx2_ASAP7_75t_R register___U10186 ( .A(Reg_data[658]), .Y(register__n6561) );
  BUFx2_ASAP7_75t_R register___U10187 ( .A(register__n10448), .Y(register__n6562) );
  BUFx4f_ASAP7_75t_R register___U10188 ( .A(register__n10448), .Y(register__n6563) );
  BUFx3_ASAP7_75t_R register___U10189 ( .A(register__n10448), .Y(register__n6564) );
  BUFx3_ASAP7_75t_R register___U10190 ( .A(register__n6566), .Y(register__n6565) );
  BUFx2_ASAP7_75t_R register___U10191 ( .A(Reg_data[648]), .Y(register__n6566) );
  BUFx3_ASAP7_75t_R register___U10192 ( .A(register__net112504), .Y(register__net112503) );
  BUFx2_ASAP7_75t_R register___U10193 ( .A(Reg_data[646]), .Y(register__net112504) );
  BUFx3_ASAP7_75t_R register___U10194 ( .A(register__net112500), .Y(register__net112499) );
  BUFx2_ASAP7_75t_R register___U10195 ( .A(Reg_data[645]), .Y(register__net112500) );
  BUFx3_ASAP7_75t_R register___U10196 ( .A(register__net112496), .Y(register__net112495) );
  BUFx2_ASAP7_75t_R register___U10197 ( .A(Reg_data[614]), .Y(register__net112496) );
  BUFx3_ASAP7_75t_R register___U10198 ( .A(register__n6568), .Y(register__n6567) );
  BUFx2_ASAP7_75t_R register___U10199 ( .A(Reg_data[611]), .Y(register__n6568) );
  BUFx3_ASAP7_75t_R register___U10200 ( .A(register__n6570), .Y(register__n6569) );
  BUFx2_ASAP7_75t_R register___U10201 ( .A(Reg_data[609]), .Y(register__n6570) );
  BUFx3_ASAP7_75t_R register___U10202 ( .A(register__n6572), .Y(register__n6571) );
  BUFx2_ASAP7_75t_R register___U10203 ( .A(Reg_data[514]), .Y(register__n6572) );
  BUFx3_ASAP7_75t_R register___U10204 ( .A(register__n6574), .Y(register__n6573) );
  BUFx2_ASAP7_75t_R register___U10205 ( .A(Reg_data[436]), .Y(register__n6574) );
  BUFx3_ASAP7_75t_R register___U10206 ( .A(register__n6576), .Y(register__n6575) );
  BUFx2_ASAP7_75t_R register___U10207 ( .A(Reg_data[434]), .Y(register__n6576) );
  BUFx3_ASAP7_75t_R register___U10208 ( .A(register__n6578), .Y(register__n6577) );
  BUFx2_ASAP7_75t_R register___U10209 ( .A(Reg_data[354]), .Y(register__n6578) );
  BUFx3_ASAP7_75t_R register___U10210 ( .A(register__n6580), .Y(register__n6579) );
  BUFx2_ASAP7_75t_R register___U10211 ( .A(Reg_data[160]), .Y(register__n6580) );
  BUFx3_ASAP7_75t_R register___U10212 ( .A(register__n6582), .Y(register__n6581) );
  BUFx2_ASAP7_75t_R register___U10213 ( .A(Reg_data[150]), .Y(register__n6582) );
  BUFx3_ASAP7_75t_R register___U10214 ( .A(register__n6584), .Y(register__n6583) );
  BUFx2_ASAP7_75t_R register___U10215 ( .A(Reg_data[148]), .Y(register__n6584) );
  BUFx3_ASAP7_75t_R register___U10216 ( .A(register__net112456), .Y(register__net112455) );
  BUFx2_ASAP7_75t_R register___U10217 ( .A(Reg_data[146]), .Y(register__net112456) );
  BUFx3_ASAP7_75t_R register___U10218 ( .A(register__n6586), .Y(register__n6585) );
  BUFx2_ASAP7_75t_R register___U10219 ( .A(Reg_data[144]), .Y(register__n6586) );
  BUFx3_ASAP7_75t_R register___U10220 ( .A(register__n6588), .Y(register__n6587) );
  BUFx2_ASAP7_75t_R register___U10221 ( .A(Reg_data[136]), .Y(register__n6588) );
  BUFx3_ASAP7_75t_R register___U10222 ( .A(register__n6590), .Y(register__n6589) );
  BUFx2_ASAP7_75t_R register___U10223 ( .A(Reg_data[129]), .Y(register__n6590) );
  BUFx3_ASAP7_75t_R register___U10224 ( .A(register__n6592), .Y(register__n6591) );
  BUFx2_ASAP7_75t_R register___U10225 ( .A(Reg_data[128]), .Y(register__n6592) );
  BUFx3_ASAP7_75t_R register___U10226 ( .A(register__n6594), .Y(register__n6593) );
  BUFx2_ASAP7_75t_R register___U10227 ( .A(Reg_data[131]), .Y(register__n6594) );
  BUFx3_ASAP7_75t_R register___U10228 ( .A(register__n6596), .Y(register__n6595) );
  BUFx2_ASAP7_75t_R register___U10229 ( .A(Reg_data[245]), .Y(register__n6596) );
  BUFx3_ASAP7_75t_R register___U10230 ( .A(register__net112428), .Y(register__net112427) );
  BUFx2_ASAP7_75t_R register___U10231 ( .A(Reg_data[632]), .Y(register__net112428) );
  BUFx3_ASAP7_75t_R register___U10232 ( .A(register__n6598), .Y(register__n6597) );
  BUFx2_ASAP7_75t_R register___U10233 ( .A(Reg_data[977]), .Y(register__n6598) );
  BUFx3_ASAP7_75t_R register___U10234 ( .A(register__net112420), .Y(register__net112419) );
  BUFx2_ASAP7_75t_R register___U10235 ( .A(Reg_data[367]), .Y(register__net112420) );
  BUFx3_ASAP7_75t_R register___U10236 ( .A(register__n6600), .Y(register__n6599) );
  BUFx2_ASAP7_75t_R register___U10237 ( .A(Reg_data[457]), .Y(register__n6600) );
  BUFx3_ASAP7_75t_R register___U10238 ( .A(register__n6602), .Y(register__n6601) );
  BUFx2_ASAP7_75t_R register___U10239 ( .A(Reg_data[620]), .Y(register__n6602) );
  BUFx3_ASAP7_75t_R register___U10240 ( .A(register__net112408), .Y(register__net112407) );
  BUFx2_ASAP7_75t_R register___U10241 ( .A(Reg_data[395]), .Y(register__net112408) );
  BUFx3_ASAP7_75t_R register___U10242 ( .A(register__n6604), .Y(register__n6603) );
  BUFx2_ASAP7_75t_R register___U10243 ( .A(Reg_data[987]), .Y(register__n6604) );
  BUFx6f_ASAP7_75t_R register___U10244 ( .A(register__n10515), .Y(register__n6606) );
  AO22x1_ASAP7_75t_R register___U10245 ( .A1(register__n6606), .A2(register__net128121), .B1(register__n8201), .B2(
        n2001), .Y(register__n11646) );
  BUFx3_ASAP7_75t_R register___U10246 ( .A(register__n6608), .Y(register__n6607) );
  BUFx2_ASAP7_75t_R register___U10247 ( .A(Reg_data[525]), .Y(register__n6608) );
  BUFx2_ASAP7_75t_R register___U10248 ( .A(register__n10130), .Y(register__n6609) );
  BUFx4f_ASAP7_75t_R register___U10249 ( .A(register__n10130), .Y(register__n6610) );
  BUFx3_ASAP7_75t_R register___U10250 ( .A(register__n6612), .Y(register__n6611) );
  BUFx2_ASAP7_75t_R register___U10251 ( .A(Reg_data[380]), .Y(register__n6612) );
  BUFx3_ASAP7_75t_R register___U10252 ( .A(register__net112382), .Y(register__net112381) );
  BUFx2_ASAP7_75t_R register___U10253 ( .A(Reg_data[618]), .Y(register__net112382) );
  BUFx3_ASAP7_75t_R register___U10254 ( .A(register__n6614), .Y(register__n6613) );
  BUFx2_ASAP7_75t_R register___U10255 ( .A(Reg_data[493]), .Y(register__n6614) );
  BUFx3_ASAP7_75t_R register___U10256 ( .A(register__n6616), .Y(register__n6615) );
  BUFx2_ASAP7_75t_R register___U10257 ( .A(Reg_data[492]), .Y(register__n6616) );
  BUFx3_ASAP7_75t_R register___U10258 ( .A(register__n6618), .Y(register__n6617) );
  BUFx2_ASAP7_75t_R register___U10259 ( .A(Reg_data[488]), .Y(register__n6618) );
  BUFx4f_ASAP7_75t_R register___U10260 ( .A(register__n9288), .Y(register__n6619) );
  BUFx2_ASAP7_75t_R register___U10261 ( .A(register__n9288), .Y(register__n6620) );
  BUFx2_ASAP7_75t_R register___U10262 ( .A(register__n9288), .Y(register__n6621) );
  BUFx3_ASAP7_75t_R register___U10263 ( .A(register__n6623), .Y(register__n6622) );
  BUFx2_ASAP7_75t_R register___U10264 ( .A(Reg_data[137]), .Y(register__n6623) );
  BUFx2_ASAP7_75t_R register___U10265 ( .A(register__n8356), .Y(register__n6624) );
  BUFx2_ASAP7_75t_R register___U10266 ( .A(register__n8356), .Y(register__n6625) );
  BUFx3_ASAP7_75t_R register___U10267 ( .A(register__net112344), .Y(register__net112343) );
  BUFx2_ASAP7_75t_R register___U10268 ( .A(Reg_data[536]), .Y(register__net112344) );
  BUFx2_ASAP7_75t_R register___U10269 ( .A(register__net89425), .Y(register__net112345) );
  BUFx4f_ASAP7_75t_R register___U10270 ( .A(register__net89425), .Y(register__net112347) );
  BUFx3_ASAP7_75t_R register___U10271 ( .A(register__net112340), .Y(register__net112339) );
  BUFx2_ASAP7_75t_R register___U10272 ( .A(Reg_data[248]), .Y(register__net112340) );
  BUFx3_ASAP7_75t_R register___U10273 ( .A(register__net112336), .Y(register__net112335) );
  BUFx2_ASAP7_75t_R register___U10274 ( .A(Reg_data[495]), .Y(register__net112336) );
  BUFx3_ASAP7_75t_R register___U10275 ( .A(register__n6628), .Y(register__n6627) );
  BUFx2_ASAP7_75t_R register___U10276 ( .A(Reg_data[135]), .Y(register__n6628) );
  BUFx2_ASAP7_75t_R register___U10277 ( .A(register__n10177), .Y(register__n6629) );
  BUFx2_ASAP7_75t_R register___U10278 ( .A(register__n10177), .Y(register__n6630) );
  BUFx4f_ASAP7_75t_R register___U10279 ( .A(register__n10177), .Y(register__n6631) );
  BUFx3_ASAP7_75t_R register___U10280 ( .A(register__n6633), .Y(register__n6632) );
  BUFx2_ASAP7_75t_R register___U10281 ( .A(Reg_data[647]), .Y(register__n6633) );
  BUFx3_ASAP7_75t_R register___U10282 ( .A(register__n6635), .Y(register__n6634) );
  BUFx2_ASAP7_75t_R register___U10283 ( .A(Reg_data[238]), .Y(register__n6635) );
  BUFx3_ASAP7_75t_R register___U10284 ( .A(register__net112314), .Y(register__net112313) );
  BUFx2_ASAP7_75t_R register___U10285 ( .A(Reg_data[221]), .Y(register__net112314) );
  BUFx3_ASAP7_75t_R register___U10286 ( .A(register__n6637), .Y(register__n6636) );
  BUFx2_ASAP7_75t_R register___U10287 ( .A(Reg_data[542]), .Y(register__n6637) );
  BUFx3_ASAP7_75t_R register___U10288 ( .A(register__n6639), .Y(register__n6638) );
  BUFx2_ASAP7_75t_R register___U10289 ( .A(Reg_data[702]), .Y(register__n6639) );
  BUFx3_ASAP7_75t_R register___U10290 ( .A(register__net112296), .Y(register__net112295) );
  BUFx2_ASAP7_75t_R register___U10291 ( .A(Reg_data[522]), .Y(register__net112296) );
  BUFx4f_ASAP7_75t_R register___U10292 ( .A(register__net89281), .Y(register__net112297) );
  BUFx2_ASAP7_75t_R register___U10293 ( .A(register__net89281), .Y(register__net112298) );
  BUFx3_ASAP7_75t_R register___U10294 ( .A(register__n6641), .Y(register__n6640) );
  BUFx2_ASAP7_75t_R register___U10295 ( .A(Reg_data[371]), .Y(register__n6641) );
  BUFx3_ASAP7_75t_R register___U10296 ( .A(register__net112282), .Y(register__net112281) );
  BUFx2_ASAP7_75t_R register___U10297 ( .A(Reg_data[490]), .Y(register__net112282) );
  BUFx4f_ASAP7_75t_R register___U10298 ( .A(register__net93456), .Y(register__net112283) );
  BUFx2_ASAP7_75t_R register___U10299 ( .A(register__net93456), .Y(register__net112285) );
  BUFx3_ASAP7_75t_R register___U10300 ( .A(register__n6643), .Y(register__n6642) );
  BUFx2_ASAP7_75t_R register___U10301 ( .A(Reg_data[151]), .Y(register__n6643) );
  BUFx2_ASAP7_75t_R register___U10302 ( .A(register__n10251), .Y(register__n6644) );
  BUFx2_ASAP7_75t_R register___U10303 ( .A(register__n10251), .Y(register__n6645) );
  BUFx4f_ASAP7_75t_R register___U10304 ( .A(register__n10251), .Y(register__n6646) );
  BUFx3_ASAP7_75t_R register___U10305 ( .A(register__n6648), .Y(register__n6647) );
  BUFx2_ASAP7_75t_R register___U10306 ( .A(Reg_data[663]), .Y(register__n6648) );
  BUFx2_ASAP7_75t_R register___U10307 ( .A(register__n10259), .Y(register__n6649) );
  BUFx2_ASAP7_75t_R register___U10308 ( .A(register__n10259), .Y(register__n6650) );
  BUFx4f_ASAP7_75t_R register___U10309 ( .A(register__n10259), .Y(register__n6651) );
  BUFx3_ASAP7_75t_R register___U10310 ( .A(register__n6653), .Y(register__n6652) );
  BUFx2_ASAP7_75t_R register___U10311 ( .A(Reg_data[503]), .Y(register__n6653) );
  BUFx3_ASAP7_75t_R register___U10312 ( .A(register__n9307), .Y(register__n6654) );
  BUFx2_ASAP7_75t_R register___U10313 ( .A(register__n9307), .Y(register__n6655) );
  BUFx4f_ASAP7_75t_R register___U10314 ( .A(register__n9307), .Y(register__n6656) );
  BUFx3_ASAP7_75t_R register___U10315 ( .A(register__n6658), .Y(register__n6657) );
  BUFx2_ASAP7_75t_R register___U10316 ( .A(Reg_data[731]), .Y(register__n6658) );
  BUFx3_ASAP7_75t_R register___U10317 ( .A(register__n6660), .Y(register__n6659) );
  BUFx2_ASAP7_75t_R register___U10318 ( .A(Reg_data[154]), .Y(register__n6660) );
  BUFx2_ASAP7_75t_R register___U10319 ( .A(register__n10279), .Y(register__n6661) );
  BUFx2_ASAP7_75t_R register___U10320 ( .A(register__n10279), .Y(register__n6662) );
  BUFx4f_ASAP7_75t_R register___U10321 ( .A(register__n10279), .Y(register__n6663) );
  BUFx3_ASAP7_75t_R register___U10322 ( .A(register__n6665), .Y(register__n6664) );
  BUFx2_ASAP7_75t_R register___U10323 ( .A(Reg_data[745]), .Y(register__n6665) );
  BUFx3_ASAP7_75t_R register___U10324 ( .A(register__n6667), .Y(register__n6666) );
  BUFx2_ASAP7_75t_R register___U10325 ( .A(Reg_data[497]), .Y(register__n6667) );
  BUFx4f_ASAP7_75t_R register___U10326 ( .A(register__n9313), .Y(register__n6668) );
  BUFx2_ASAP7_75t_R register___U10327 ( .A(register__n9313), .Y(register__n6669) );
  BUFx2_ASAP7_75t_R register___U10328 ( .A(register__n9313), .Y(register__n6670) );
  BUFx3_ASAP7_75t_R register___U10329 ( .A(register__n6672), .Y(register__n6671) );
  BUFx2_ASAP7_75t_R register___U10330 ( .A(Reg_data[507]), .Y(register__n6672) );
  BUFx3_ASAP7_75t_R register___U10331 ( .A(register__n6674), .Y(register__n6673) );
  BUFx2_ASAP7_75t_R register___U10332 ( .A(Reg_data[63]), .Y(register__n6674) );
  BUFx3_ASAP7_75t_R register___U10333 ( .A(register__n6676), .Y(register__n6675) );
  BUFx2_ASAP7_75t_R register___U10334 ( .A(Reg_data[255]), .Y(register__n6676) );
  BUFx3_ASAP7_75t_R register___U10335 ( .A(register__net112208), .Y(register__net112207) );
  BUFx2_ASAP7_75t_R register___U10336 ( .A(Reg_data[61]), .Y(register__net112208) );
  BUFx3_ASAP7_75t_R register___U10337 ( .A(register__n6678), .Y(register__n6677) );
  BUFx2_ASAP7_75t_R register___U10338 ( .A(Reg_data[398]), .Y(register__n6678) );
  BUFx4f_ASAP7_75t_R register___U10339 ( .A(register__net97245), .Y(register__C6423_net60596) );
  INVx1_ASAP7_75t_R register___U10340 ( .A(register__C6423_net60596), .Y(register__net112155) );
  BUFx6f_ASAP7_75t_R register___U10341 ( .A(register__net97246), .Y(register__net97245) );
  BUFx4f_ASAP7_75t_R register___U10342 ( .A(register__n3447), .Y(register__n12299) );
  BUFx6f_ASAP7_75t_R register___U10343 ( .A(register__n6680), .Y(register__n12137) );
  BUFx6f_ASAP7_75t_R register___U10344 ( .A(register__n6680), .Y(register__n12139) );
  BUFx4f_ASAP7_75t_R register___U10345 ( .A(register__n6680), .Y(register__n12140) );
  OA22x2_ASAP7_75t_R register___U10346 ( .A1(register__net63258), .A2(register__n110), .B1(register__net88785), .B2(
        n1665), .Y(register__n12640) );
  OA22x2_ASAP7_75t_R register___U10347 ( .A1(register__n12063), .A2(register__n7327), .B1(register__n9587), .B2(register__n12504), 
        .Y(register__n12570) );
  OA22x2_ASAP7_75t_R register___U10348 ( .A1(register__n12052), .A2(register__n1709), .B1(register__n10008), .B2(register__n3353), 
        .Y(register__n13256) );
  INVx1_ASAP7_75t_R register___U10349 ( .A(register__n4872), .Y(register__n6681) );
  OA22x2_ASAP7_75t_R register___U10350 ( .A1(register__n11950), .A2(register__n399), .B1(register__n10454), .B2(register__n11742), 
        .Y(register__n13305) );
  OA22x2_ASAP7_75t_R register___U10351 ( .A1(register__n12151), .A2(register__n7327), .B1(register__n9754), .B2(register__n3540), 
        .Y(register__n12566) );
  INVx1_ASAP7_75t_R register___U10352 ( .A(register__n12566), .Y(register__n6684) );
  OA22x2_ASAP7_75t_R register___U10353 ( .A1(register__n12144), .A2(register__n1738), .B1(register__n10148), .B2(register__n3681), 
        .Y(register__n13251) );
  OA22x2_ASAP7_75t_R register___U10354 ( .A1(register__net64020), .A2(register__n7327), .B1(register__net90529), .B2(
        n7973), .Y(register__n12564) );
  OA22x2_ASAP7_75t_R register___U10355 ( .A1(register__net63996), .A2(register__n1720), .B1(register__net89405), .B2(
        n11870), .Y(register__n13250) );
  OA22x2_ASAP7_75t_R register___U10356 ( .A1(register__n12396), .A2(register__n1707), .B1(register__n10281), .B2(register__n1719), 
        .Y(register__n13243) );
  OA22x2_ASAP7_75t_R register___U10357 ( .A1(register__net62652), .A2(register__n1725), .B1(register__n10295), .B2(
        n1692), .Y(register__n13239) );
  OA22x2_ASAP7_75t_R register___U10358 ( .A1(register__n12395), .A2(register__n399), .B1(register__n10303), .B2(register__n8334), 
        .Y(register__n13290) );
  OA22x2_ASAP7_75t_R register___U10359 ( .A1(register__net63256), .A2(register__n665), .B1(register__net89045), .B2(register__n81), .Y(register__n12807) );
  INVx1_ASAP7_75t_R register___U10360 ( .A(register__n5405), .Y(register__n6687) );
  OA22x2_ASAP7_75t_R register___U10361 ( .A1(register__n12430), .A2(register__n2801), .B1(register__n10335), .B2(register__n3076), 
        .Y(register__n12803) );
  OA22x2_ASAP7_75t_R register___U10362 ( .A1(register__n12233), .A2(register__n665), .B1(register__n10313), .B2(register__n81), 
        .Y(register__n12814) );
  OA22x2_ASAP7_75t_R register___U10363 ( .A1(register__n12430), .A2(register__n4033), .B1(register__n9345), .B2(register__n3359), 
        .Y(register__n12525) );
  OA22x2_ASAP7_75t_R register___U10364 ( .A1(register__net64354), .A2(register__n117), .B1(register__net106199), .B2(
        n1671), .Y(register__n12652) );
  INVx1_ASAP7_75t_R register___U10365 ( .A(register__n4405), .Y(register__n6690) );
  OA22x2_ASAP7_75t_R register___U10366 ( .A1(register__n12426), .A2(register__n894), .B1(register__n7522), .B2(register__n907), 
        .Y(register__n13040) );
  INVx1_ASAP7_75t_R register___U10367 ( .A(register__n13040), .Y(register__n6691) );
  OA22x2_ASAP7_75t_R register___U10368 ( .A1(register__net64424), .A2(register__n891), .B1(register__net101004), .B2(
        n901), .Y(register__n13055) );
  OA22x2_ASAP7_75t_R register___U10369 ( .A1(register__n12407), .A2(register__n119), .B1(register__n8516), .B2(register__n1536), 
        .Y(register__n12583) );
  OA22x2_ASAP7_75t_R register___U10370 ( .A1(register__net62658), .A2(register__n1092), .B1(register__n7574), .B2(register__n3675), .Y(register__n13064) );
  INVx1_ASAP7_75t_R register___U10371 ( .A(register__n4892), .Y(register__n6693) );
  OA22x2_ASAP7_75t_R register___U10372 ( .A1(register__net64328), .A2(register__n1092), .B1(register__net90669), .B2(
        n5531), .Y(register__n13080) );
  OA22x2_ASAP7_75t_R register___U10373 ( .A1(register__n12081), .A2(register__n399), .B1(register__n10275), .B2(register__n12486), 
        .Y(register__n13301) );
  INVx1_ASAP7_75t_R register___U10374 ( .A(register__n4888), .Y(register__n6694) );
  OA22x2_ASAP7_75t_R register___U10375 ( .A1(register__net62844), .A2(register__n7327), .B1(register__net90213), .B2(
        n11836), .Y(register__n12555) );
  INVx1_ASAP7_75t_R register___U10376 ( .A(register__n4599), .Y(register__n6695) );
  OA22x2_ASAP7_75t_R register___U10377 ( .A1(register__n12421), .A2(register__n399), .B1(register__n10223), .B2(register__n1161), 
        .Y(register__n13288) );
  INVx1_ASAP7_75t_R register___U10378 ( .A(register__n5609), .Y(register__n6698) );
  INVx1_ASAP7_75t_R register___U10379 ( .A(register__n5801), .Y(register__n6700) );
  INVx1_ASAP7_75t_R register___U10380 ( .A(register__n4447), .Y(register__n6703) );
  INVx1_ASAP7_75t_R register___U10381 ( .A(register__n4449), .Y(register__n6704) );
  INVx1_ASAP7_75t_R register___U10382 ( .A(register__n4807), .Y(register__n6706) );
  INVx1_ASAP7_75t_R register___U10383 ( .A(register__n4809), .Y(register__n6707) );
  INVx1_ASAP7_75t_R register___U10384 ( .A(register__n5601), .Y(register__n6708) );
  INVx1_ASAP7_75t_R register___U10385 ( .A(register__n5603), .Y(register__n6710) );
  INVx1_ASAP7_75t_R register___U10386 ( .A(register__n4718), .Y(register__n6712) );
  INVx1_ASAP7_75t_R register___U10387 ( .A(register__n5584), .Y(register__n6714) );
  INVx1_ASAP7_75t_R register___U10388 ( .A(register__n10566), .Y(register__n6715) );
  INVx1_ASAP7_75t_R register___U10389 ( .A(register__n4793), .Y(register__n6716) );
  INVx1_ASAP7_75t_R register___U10390 ( .A(register__n10771), .Y(register__n6718) );
  BUFx12f_ASAP7_75t_R register___U10391 ( .A(register__n4841), .Y(register__n11824) );
  BUFx12f_ASAP7_75t_R register___U10392 ( .A(register__n5182), .Y(register__n11850) );
  BUFx12f_ASAP7_75t_R register___U10393 ( .A(register__n4373), .Y(register__n11733) );
  OA22x2_ASAP7_75t_R register___U10394 ( .A1(register__n12349), .A2(register__n7327), .B1(register__n7399), .B2(register__n11914), 
        .Y(register__n12560) );
  INVx1_ASAP7_75t_R register___U10395 ( .A(register__n5958), .Y(register__n6722) );
  OA22x2_ASAP7_75t_R register___U10396 ( .A1(register__net64356), .A2(register__n119), .B1(register__net95342), .B2(
        n1538), .Y(register__n12596) );
  OA22x2_ASAP7_75t_R register___U10397 ( .A1(register__n12056), .A2(register__n891), .B1(register__n10493), .B2(register__n906), 
        .Y(register__n13057) );
  INVx1_ASAP7_75t_R register___U10398 ( .A(register__n5755), .Y(register__n6723) );
  OA22x2_ASAP7_75t_R register___U10399 ( .A1(register__n12323), .A2(register__n107), .B1(register__n8343), .B2(register__n1519), 
        .Y(register__n12588) );
  OA22x2_ASAP7_75t_R register___U10400 ( .A1(register__n12262), .A2(register__n11829), .B1(register__net91045), .B2(
        n1523), .Y(register__n12590) );
  INVx1_ASAP7_75t_R register___U10401 ( .A(register__n3853), .Y(register__n6725) );
  OA22x2_ASAP7_75t_R register___U10402 ( .A1(register__n12063), .A2(register__n2008), .B1(register__n9601), .B2(register__n1531), 
        .Y(register__n12598) );
  OA22x2_ASAP7_75t_R register___U10403 ( .A1(register__n11959), .A2(register__n1946), .B1(register__n9359), .B2(register__n3746), 
        .Y(register__n12830) );
  OA22x2_ASAP7_75t_R register___U10404 ( .A1(register__n12316), .A2(register__n894), .B1(register__n9662), .B2(register__n897), 
        .Y(register__n13046) );
  OA22x2_ASAP7_75t_R register___U10405 ( .A1(register__n11989), .A2(register__n893), .B1(register__n9666), .B2(register__n906), 
        .Y(register__n13062) );
  OA22x2_ASAP7_75t_R register___U10406 ( .A1(register__n12236), .A2(register__n1548), .B1(register__n7992), .B2(register__n1543), 
        .Y(register__n12591) );
  OA22x2_ASAP7_75t_R register___U10407 ( .A1(register__n3759), .A2(register__n4033), .B1(register__n9573), .B2(register__n11839), 
        .Y(register__n12537) );
  INVx1_ASAP7_75t_R register___U10408 ( .A(register__n3757), .Y(register__n6730) );
  OA22x2_ASAP7_75t_R register___U10409 ( .A1(register__net64776), .A2(register__n107), .B1(register__net91033), .B2(
        n1526), .Y(register__n12600) );
  OA22x2_ASAP7_75t_R register___U10410 ( .A1(register__n12031), .A2(register__n1549), .B1(register__n9603), .B2(register__n1535), 
        .Y(register__n12603) );
  OA22x2_ASAP7_75t_R register___U10411 ( .A1(register__register__n11934), .A2(register__n119), .B1(register__n9605), .B2(register__n1539), 
        .Y(register__n12605) );
  OA22x2_ASAP7_75t_R register___U10412 ( .A1(register__n11962), .A2(register__n111), .B1(register__n8330), .B2(register__n1672), 
        .Y(register__n12659) );
  OA22x2_ASAP7_75t_R register___U10413 ( .A1(register__net64940), .A2(register__n1991), .B1(register__n9209), .B2(register__n1602), .Y(register__n12713) );
  OA22x2_ASAP7_75t_R register___U10414 ( .A1(register__net64928), .A2(register__n893), .B1(register__n9664), .B2(register__n902), 
        .Y(register__n13060) );
  INVx1_ASAP7_75t_R register___U10415 ( .A(register__n5083), .Y(register__n6733) );
  OA22x2_ASAP7_75t_R register___U10416 ( .A1(register__net64674), .A2(register__n1092), .B1(register__n9726), .B2(register__n3511), .Y(register__n13082) );
  INVx1_ASAP7_75t_R register___U10417 ( .A(register__n4214), .Y(register__n6734) );
  OA22x2_ASAP7_75t_R register___U10418 ( .A1(register__net63266), .A2(register__n4033), .B1(register__net93793), .B2(
        n3736), .Y(register__n12529) );
  INVx1_ASAP7_75t_R register___U10419 ( .A(register__n6242), .Y(register__n6735) );
  OA22x2_ASAP7_75t_R register___U10420 ( .A1(register__net63254), .A2(register__n2815), .B1(register__net91335), .B2(
        n1925), .Y(register__n12865) );
  INVx1_ASAP7_75t_R register___U10421 ( .A(register__n6244), .Y(register__n6736) );
  OA22x2_ASAP7_75t_R register___U10422 ( .A1(register__net64436), .A2(register__n3022), .B1(register__net97177), .B2(
        n884), .Y(register__n12708) );
  INVx4_ASAP7_75t_R register___U10423 ( .A(register__net64472), .Y(register__net64436) );
  OA22x2_ASAP7_75t_R register___U10424 ( .A1(register__net64018), .A2(register__n114), .B1(register__net91307), .B2(
        n1668), .Y(register__n12648) );
  OA22x2_ASAP7_75t_R register___U10425 ( .A1(register__n12119), .A2(register__n1927), .B1(register__n9529), .B2(register__n1939), 
        .Y(register__n12876) );
  INVx1_ASAP7_75t_R register___U10426 ( .A(register__n5576), .Y(register__n6738) );
  OA22x2_ASAP7_75t_R register___U10427 ( .A1(register__net63344), .A2(register__n3022), .B1(register__n9533), .B2(register__n1589), .Y(register__n12697) );
  INVx1_ASAP7_75t_R register___U10428 ( .A(register__n4669), .Y(register__n6739) );
  OA22x2_ASAP7_75t_R register___U10429 ( .A1(register__n12402), .A2(register__n1942), .B1(register__n9537), .B2(register__n1937), 
        .Y(register__n12863) );
  OA22x2_ASAP7_75t_R register___U10430 ( .A1(register__n12285), .A2(register__n892), .B1(register__n9760), .B2(register__n903), 
        .Y(register__n13047) );
  INVx2_ASAP7_75t_R register___U10431 ( .A(register__n12299), .Y(register__n12285) );
  OA22x2_ASAP7_75t_R register___U10432 ( .A1(register__net124970), .A2(register__n892), .B1(register__n8811), .B2(register__n905), 
        .Y(register__n13041) );
  OA22x2_ASAP7_75t_R register___U10433 ( .A1(register__n12092), .A2(register__n117), .B1(register__n7997), .B2(register__n1660), 
        .Y(register__n12654) );
  INVx1_ASAP7_75t_R register___U10434 ( .A(register__n5089), .Y(register__n6742) );
  INVx3_ASAP7_75t_R register___U10435 ( .A(register__net64724), .Y(register__net64690) );
  OA22x2_ASAP7_75t_R register___U10436 ( .A1(register__net64432), .A2(register__n1069), .B1(register__net89277), .B2(
        n81), .Y(register__n12821) );
  INVx1_ASAP7_75t_R register___U10437 ( .A(register__n3777), .Y(register__n6743) );
  OA22x2_ASAP7_75t_R register___U10438 ( .A1(register__n12403), .A2(register__n1069), .B1(register__n10287), .B2(register__n3076), 
        .Y(register__n12805) );
  OA22x2_ASAP7_75t_R register___U10439 ( .A1(register__net62834), .A2(register__n2819), .B1(register__net94144), .B2(
        n1928), .Y(register__n12861) );
  OA22x2_ASAP7_75t_R register___U10440 ( .A1(register__net109773), .A2(register__n665), .B1(register__n4962), .B2(register__n3076), .Y(register__n12800) );
  INVx1_ASAP7_75t_R register___U10441 ( .A(register__n4221), .Y(register__n6745) );
  INVx1_ASAP7_75t_R register___U10442 ( .A(register__n4223), .Y(register__n6746) );
  INVx1_ASAP7_75t_R register___U10443 ( .A(register__n4721), .Y(register__n6748) );
  AO22x1_ASAP7_75t_R register___U10444 ( .A1(register__n10479), .A2(register__C6423_net61318), .B1(register__n10452), 
        .B2(register__C6423_net72545), .Y(register__n11551) );
  INVx1_ASAP7_75t_R register___U10445 ( .A(register__n4580), .Y(register__n6749) );
  INVx1_ASAP7_75t_R register___U10446 ( .A(register__n4050), .Y(register__n6750) );
  OA22x2_ASAP7_75t_R register___U10447 ( .A1(register__n3665), .A2(register__n110), .B1(register__n9441), .B2(register__n1678), 
        .Y(register__n12657) );
  OA22x2_ASAP7_75t_R register___U10448 ( .A1(register__n4045), .A2(register__n2935), .B1(register__n9453), .B2(register__n1596), 
        .Y(register__n12714) );
  INVx1_ASAP7_75t_R register___U10449 ( .A(register__n4651), .Y(register__n6755) );
  OA22x2_ASAP7_75t_R register___U10450 ( .A1(register__n4999), .A2(register__n1957), .B1(register__n9461), .B2(register__n2807), 
        .Y(register__n12868) );
  OA22x2_ASAP7_75t_R register___U10451 ( .A1(register__net64766), .A2(register__n1921), .B1(register__net91463), .B2(
        n11884), .Y(register__n12881) );
  OA22x2_ASAP7_75t_R register___U10452 ( .A1(register__n12027), .A2(register__n2804), .B1(register__n9467), .B2(register__n1945), 
        .Y(register__n12884) );
  INVx1_ASAP7_75t_R register___U10453 ( .A(register__n5568), .Y(register__n6756) );
  BUFx12f_ASAP7_75t_R register___U10454 ( .A(register__n11738), .Y(register__n11737) );
  BUFx2_ASAP7_75t_R register___U10455 ( .A(register__n11227), .Y(register__n6762) );
  INVx2_ASAP7_75t_R register___U10456 ( .A(register__n7780), .Y(register__n6764) );
  BUFx2_ASAP7_75t_R register___U10457 ( .A(register__n10531), .Y(register__n6765) );
  BUFx2_ASAP7_75t_R register___U10458 ( .A(register__n10596), .Y(register__n6766) );
  INVx2_ASAP7_75t_R register___U10459 ( .A(register__n9477), .Y(register__n10936) );
  BUFx2_ASAP7_75t_R register___U10460 ( .A(register__n11524), .Y(register__n6767) );
  BUFx2_ASAP7_75t_R register___U10461 ( .A(register__n11479), .Y(register__n6768) );
  BUFx2_ASAP7_75t_R register___U10462 ( .A(register__n11202), .Y(register__n6769) );
  BUFx2_ASAP7_75t_R register___U10463 ( .A(register__n11160), .Y(register__n6770) );
  BUFx2_ASAP7_75t_R register___U10464 ( .A(register__n10933), .Y(register__n6771) );
  INVx2_ASAP7_75t_R register___U10465 ( .A(register__n9463), .Y(register__n11525) );
  BUFx2_ASAP7_75t_R register___U10466 ( .A(register__n10867), .Y(register__n6772) );
  BUFx2_ASAP7_75t_R register___U10467 ( .A(register__C6422_net59855), .Y(register__net111143) );
  BUFx2_ASAP7_75t_R register___U10468 ( .A(register__n10761), .Y(register__n6773) );
  INVx2_ASAP7_75t_R register___U10469 ( .A(register__n10387), .Y(register__n11686) );
  INVx2_ASAP7_75t_R register___U10470 ( .A(register__n9531), .Y(register__n11501) );
  INVx2_ASAP7_75t_R register___U10471 ( .A(register__n10383), .Y(register__n11061) );
  BUFx2_ASAP7_75t_R register___U10472 ( .A(register__C6423_net61113), .Y(register__net111131) );
  INVx2_ASAP7_75t_R register___U10473 ( .A(register__n9563), .Y(register__n10890) );
  INVx2_ASAP7_75t_R register___U10474 ( .A(register__n9525), .Y(register__n11104) );
  INVx2_ASAP7_75t_R register___U10475 ( .A(register__n9535), .Y(register__n11644) );
  BUFx2_ASAP7_75t_R register___U10476 ( .A(register__n11583), .Y(register__n6774) );
  BUFx4f_ASAP7_75t_R register___U10477 ( .A(register__n8588), .Y(register__n6775) );
  BUFx2_ASAP7_75t_R register___U10478 ( .A(register__n8588), .Y(register__n6776) );
  BUFx2_ASAP7_75t_R register___U10479 ( .A(register__n8588), .Y(register__n6777) );
  INVx1_ASAP7_75t_R register___U10480 ( .A(register__n10415), .Y(register__n11126) );
  BUFx2_ASAP7_75t_R register___U10481 ( .A(register__n6784), .Y(register__n6783) );
  BUFx2_ASAP7_75t_R register___U10482 ( .A(register__n6788), .Y(register__n6787) );
  BUFx2_ASAP7_75t_R register___U10483 ( .A(register__n12682), .Y(register__n6788) );
  BUFx2_ASAP7_75t_R register___U10484 ( .A(register__n6792), .Y(register__n6791) );
  BUFx2_ASAP7_75t_R register___U10485 ( .A(register__n13092), .Y(register__n6792) );
  BUFx2_ASAP7_75t_R register___U10486 ( .A(register__n6794), .Y(register__n6793) );
  BUFx2_ASAP7_75t_R register___U10487 ( .A(register__n13182), .Y(register__n6794) );
  BUFx2_ASAP7_75t_R register___U10488 ( .A(register__n6798), .Y(register__n6797) );
  BUFx2_ASAP7_75t_R register___U10489 ( .A(register__n13240), .Y(register__n6798) );
  BUFx2_ASAP7_75t_R register___U10490 ( .A(register__n6800), .Y(register__n6799) );
  BUFx2_ASAP7_75t_R register___U10491 ( .A(register__n13081), .Y(register__n6800) );
  OR2x2_ASAP7_75t_R register___U10492 ( .A(register__n6802), .B(register__n6803), .Y(register__n6801) );
  BUFx2_ASAP7_75t_R register___U10493 ( .A(register__n8606), .Y(register__n6802) );
  BUFx6f_ASAP7_75t_R register___U10494 ( .A(register__n7328), .Y(register__n10824) );
  BUFx6f_ASAP7_75t_R register___U10495 ( .A(register__n7330), .Y(register__n11349) );
  BUFx6f_ASAP7_75t_R register___U10496 ( .A(register__n7332), .Y(register__n10740) );
  BUFx6f_ASAP7_75t_R register___U10497 ( .A(register__n7334), .Y(register__n11623) );
  BUFx2_ASAP7_75t_R register___U10498 ( .A(Reg_data[852]), .Y(register__n6807) );
  BUFx6f_ASAP7_75t_R register___U10499 ( .A(register__n7955), .Y(register__n7954) );
  BUFx4f_ASAP7_75t_R register___U10500 ( .A(register__n6806), .Y(register__n7955) );
  BUFx3_ASAP7_75t_R register___U10501 ( .A(register__n7737), .Y(register__n6808) );
  BUFx4f_ASAP7_75t_R register___U10502 ( .A(register__net98859), .Y(register__net94169) );
  BUFx3_ASAP7_75t_R register___U10503 ( .A(register__n7386), .Y(register__n6809) );
  BUFx4f_ASAP7_75t_R register___U10504 ( .A(register__n6809), .Y(register__n8723) );
  BUFx3_ASAP7_75t_R register___U10505 ( .A(register__n7138), .Y(register__n6810) );
  BUFx3_ASAP7_75t_R register___U10506 ( .A(register__n8841), .Y(register__n6811) );
  BUFx3_ASAP7_75t_R register___U10507 ( .A(register__n9072), .Y(register__n6812) );
  BUFx4f_ASAP7_75t_R register___U10508 ( .A(register__n8380), .Y(register__n9214) );
  BUFx3_ASAP7_75t_R register___U10509 ( .A(register__n6814), .Y(register__n6813) );
  BUFx2_ASAP7_75t_R register___U10510 ( .A(Reg_data[853]), .Y(register__n6814) );
  BUFx4f_ASAP7_75t_R register___U10511 ( .A(register__n6813), .Y(register__n7983) );
  BUFx3_ASAP7_75t_R register___U10512 ( .A(register__n6816), .Y(register__n6815) );
  BUFx2_ASAP7_75t_R register___U10513 ( .A(Reg_data[850]), .Y(register__n6816) );
  BUFx4f_ASAP7_75t_R register___U10514 ( .A(register__n6815), .Y(register__n7985) );
  BUFx3_ASAP7_75t_R register___U10515 ( .A(register__n6818), .Y(register__n6817) );
  BUFx2_ASAP7_75t_R register___U10516 ( .A(Reg_data[273]), .Y(register__n6818) );
  BUFx4f_ASAP7_75t_R register___U10517 ( .A(register__n6817), .Y(register__n7662) );
  BUFx3_ASAP7_75t_R register___U10518 ( .A(register__n6820), .Y(register__n6819) );
  BUFx2_ASAP7_75t_R register___U10519 ( .A(Reg_data[270]), .Y(register__n6820) );
  BUFx4f_ASAP7_75t_R register___U10520 ( .A(register__n6819), .Y(register__n8729) );
  BUFx3_ASAP7_75t_R register___U10521 ( .A(register__n6822), .Y(register__n6821) );
  BUFx2_ASAP7_75t_R register___U10522 ( .A(Reg_data[346]), .Y(register__n6822) );
  BUFx4f_ASAP7_75t_R register___U10523 ( .A(register__n8738), .Y(register__n6823) );
  BUFx4f_ASAP7_75t_R register___U10524 ( .A(register__n8738), .Y(register__n6824) );
  BUFx4f_ASAP7_75t_R register___U10525 ( .A(register__n6821), .Y(register__n8739) );
  BUFx3_ASAP7_75t_R register___U10526 ( .A(register__net110419), .Y(register__net110418) );
  BUFx2_ASAP7_75t_R register___U10527 ( .A(Reg_data[792]), .Y(register__net110419) );
  BUFx4f_ASAP7_75t_R register___U10528 ( .A(register__net110418), .Y(register__net102360) );
  INVx1_ASAP7_75t_R register___U10529 ( .A(register__n5266), .Y(register__n6825) );
  INVx1_ASAP7_75t_R register___U10530 ( .A(register__n5070), .Y(register__n6827) );
  BUFx6f_ASAP7_75t_R register___U10531 ( .A(register__net66310), .Y(register__net66314) );
  BUFx12f_ASAP7_75t_R register___U10532 ( .A(register__net115025), .Y(register__net66310) );
  BUFx3_ASAP7_75t_R register___U10533 ( .A(register__n6832), .Y(register__n6831) );
  BUFx2_ASAP7_75t_R register___U10534 ( .A(Reg_data[981]), .Y(register__n6832) );
  BUFx3_ASAP7_75t_R register___U10535 ( .A(register__n6834), .Y(register__n6833) );
  BUFx2_ASAP7_75t_R register___U10536 ( .A(Reg_data[976]), .Y(register__n6834) );
  BUFx4f_ASAP7_75t_R register___U10537 ( .A(register__net112748), .Y(register__net110254) );
  BUFx2_ASAP7_75t_R register___U10538 ( .A(Reg_data[825]), .Y(register__net110255) );
  BUFx6f_ASAP7_75t_R register___U10539 ( .A(register__net110254), .Y(register__net91021) );
  BUFx3_ASAP7_75t_R register___U10540 ( .A(register__n6836), .Y(register__n6835) );
  BUFx2_ASAP7_75t_R register___U10541 ( .A(Reg_data[822]), .Y(register__n6836) );
  BUFx3_ASAP7_75t_R register___U10542 ( .A(register__n9607), .Y(register__n6837) );
  BUFx2_ASAP7_75t_R register___U10543 ( .A(register__n9607), .Y(register__n6838) );
  BUFx4f_ASAP7_75t_R register___U10544 ( .A(register__n9607), .Y(register__n6839) );
  BUFx3_ASAP7_75t_R register___U10545 ( .A(register__n6841), .Y(register__n6840) );
  BUFx2_ASAP7_75t_R register___U10546 ( .A(Reg_data[821]), .Y(register__n6841) );
  BUFx4f_ASAP7_75t_R register___U10547 ( .A(register__n6036), .Y(register__n6842) );
  BUFx2_ASAP7_75t_R register___U10548 ( .A(Reg_data[818]), .Y(register__n6843) );
  BUFx12f_ASAP7_75t_R register___U10549 ( .A(register__n9614), .Y(register__n9613) );
  BUFx6f_ASAP7_75t_R register___U10550 ( .A(register__n6842), .Y(register__n9614) );
  BUFx3_ASAP7_75t_R register___U10551 ( .A(register__n6845), .Y(register__n6844) );
  BUFx2_ASAP7_75t_R register___U10552 ( .A(Reg_data[739]), .Y(register__n6845) );
  BUFx3_ASAP7_75t_R register___U10553 ( .A(register__n6847), .Y(register__n6846) );
  BUFx2_ASAP7_75t_R register___U10554 ( .A(Reg_data[737]), .Y(register__n6847) );
  BUFx3_ASAP7_75t_R register___U10555 ( .A(register__n10430), .Y(register__n6848) );
  BUFx2_ASAP7_75t_R register___U10556 ( .A(register__n10430), .Y(register__n6849) );
  BUFx4f_ASAP7_75t_R register___U10557 ( .A(register__n10430), .Y(register__n6850) );
  BUFx3_ASAP7_75t_R register___U10558 ( .A(register__n6852), .Y(register__n6851) );
  BUFx2_ASAP7_75t_R register___U10559 ( .A(Reg_data[708]), .Y(register__n6852) );
  BUFx3_ASAP7_75t_R register___U10560 ( .A(register__n6854), .Y(register__n6853) );
    BUFx2_ASAP7_75t_R register___U10561 ( .A(Reg_data[640]), .Y(register__n6854) );
  BUFx12f_ASAP7_75t_R register___U10562 ( .A(register__n9952), .Y(register__n6855) );
  BUFx12f_ASAP7_75t_R register___U10563 ( .A(register__n6855), .Y(register__n9951) );
  BUFx3_ASAP7_75t_R register___U10564 ( .A(register__net110206), .Y(register__net110205) );
  BUFx2_ASAP7_75t_R register___U10565 ( .A(Reg_data[613]), .Y(register__net110206) );
  BUFx3_ASAP7_75t_R register___U10566 ( .A(register__n6857), .Y(register__n6856) );
  BUFx2_ASAP7_75t_R register___U10567 ( .A(Reg_data[608]), .Y(register__n6857) );
  BUFx3_ASAP7_75t_R register___U10568 ( .A(register__net110198), .Y(register__net110197) );
  BUFx2_ASAP7_75t_R register___U10569 ( .A(Reg_data[537]), .Y(register__net110198) );
  BUFx3_ASAP7_75t_R register___U10570 ( .A(register__n6859), .Y(register__n6858) );
  BUFx2_ASAP7_75t_R register___U10571 ( .A(Reg_data[450]), .Y(register__n6859) );
  BUFx3_ASAP7_75t_R register___U10572 ( .A(register__n6861), .Y(register__n6860) );
  BUFx2_ASAP7_75t_R register___U10573 ( .A(Reg_data[406]), .Y(register__n6861) );
  BUFx3_ASAP7_75t_R register___U10574 ( .A(register__n6863), .Y(register__n6862) );
  BUFx2_ASAP7_75t_R register___U10575 ( .A(Reg_data[392]), .Y(register__n6863) );
  BUFx3_ASAP7_75t_R register___U10576 ( .A(register__n6865), .Y(register__n6864) );
  BUFx2_ASAP7_75t_R register___U10577 ( .A(Reg_data[355]), .Y(register__n6865) );
  BUFx3_ASAP7_75t_R register___U10578 ( .A(register__n6867), .Y(register__n6866) );
  BUFx2_ASAP7_75t_R register___U10579 ( .A(Reg_data[353]), .Y(register__n6867) );
  BUFx3_ASAP7_75t_R register___U10580 ( .A(register__n6869), .Y(register__n6868) );
  BUFx2_ASAP7_75t_R register___U10581 ( .A(Reg_data[176]), .Y(register__n6869) );
  BUFx3_ASAP7_75t_R register___U10582 ( .A(register__n6871), .Y(register__n6870) );
  BUFx2_ASAP7_75t_R register___U10583 ( .A(Reg_data[72]), .Y(register__n6871) );
  BUFx3_ASAP7_75t_R register___U10584 ( .A(register__n6873), .Y(register__n6872) );
  BUFx2_ASAP7_75t_R register___U10585 ( .A(Reg_data[967]), .Y(register__n6873) );
  BUFx3_ASAP7_75t_R register___U10586 ( .A(register__n6875), .Y(register__n6874) );
  BUFx2_ASAP7_75t_R register___U10587 ( .A(Reg_data[622]), .Y(register__n6875) );
  BUFx3_ASAP7_75t_R register___U10588 ( .A(register__n10106), .Y(register__n6876) );
  BUFx4f_ASAP7_75t_R register___U10589 ( .A(register__n10106), .Y(register__n6877) );
  BUFx2_ASAP7_75t_R register___U10590 ( .A(register__n10106), .Y(register__n6878) );
  BUFx3_ASAP7_75t_R register___U10591 ( .A(register__n6880), .Y(register__n6879) );
  BUFx2_ASAP7_75t_R register___U10592 ( .A(Reg_data[77]), .Y(register__n6880) );
  BUFx3_ASAP7_75t_R register___U10593 ( .A(register__n6882), .Y(register__n6881) );
  BUFx2_ASAP7_75t_R register___U10594 ( .A(Reg_data[62]), .Y(register__n6882) );
  BUFx3_ASAP7_75t_R register___U10595 ( .A(register__n6884), .Y(register__n6883) );
  BUFx2_ASAP7_75t_R register___U10596 ( .A(Reg_data[988]), .Y(register__n6884) );
  BUFx12f_ASAP7_75t_R register___U10597 ( .A(register__n9346), .Y(register__n6885) );
  BUFx12f_ASAP7_75t_R register___U10598 ( .A(register__n6885), .Y(register__n9345) );
  BUFx3_ASAP7_75t_R register___U10599 ( .A(register__n6887), .Y(register__n6886) );
  BUFx2_ASAP7_75t_R register___U10600 ( .A(Reg_data[986]), .Y(register__n6887) );
  BUFx3_ASAP7_75t_R register___U10601 ( .A(register__n6889), .Y(register__n6888) );
  BUFx2_ASAP7_75t_R register___U10602 ( .A(Reg_data[44]), .Y(register__n6889) );
  BUFx3_ASAP7_75t_R register___U10603 ( .A(register__net110123), .Y(register__net110122) );
  BUFx2_ASAP7_75t_R register___U10604 ( .A(Reg_data[505]), .Y(register__net110123) );
  BUFx4f_ASAP7_75t_R register___U10605 ( .A(register__net93464), .Y(register__net110124) );
  BUFx2_ASAP7_75t_R register___U10606 ( .A(register__net93464), .Y(register__net110126) );
  BUFx3_ASAP7_75t_R register___U10607 ( .A(register__n6891), .Y(register__n6890) );
  BUFx2_ASAP7_75t_R register___U10608 ( .A(Reg_data[496]), .Y(register__n6891) );
  BUFx2_ASAP7_75t_R register___U10609 ( .A(register__n8773), .Y(register__n6892) );
  BUFx6f_ASAP7_75t_R register___U10610 ( .A(register__n8773), .Y(register__n6893) );
  BUFx3_ASAP7_75t_R register___U10611 ( .A(register__n6895), .Y(register__n6894) );
  BUFx2_ASAP7_75t_R register___U10612 ( .A(Reg_data[502]), .Y(register__n6895) );
  BUFx4f_ASAP7_75t_R register___U10613 ( .A(register__n9276), .Y(register__n6896) );
  BUFx2_ASAP7_75t_R register___U10614 ( .A(register__n9276), .Y(register__n6897) );
  BUFx2_ASAP7_75t_R register___U10615 ( .A(register__n9276), .Y(register__n6898) );
  BUFx3_ASAP7_75t_R register___U10616 ( .A(register__n6900), .Y(register__n6899) );
  BUFx2_ASAP7_75t_R register___U10617 ( .A(Reg_data[500]), .Y(register__n6900) );
  BUFx3_ASAP7_75t_R register___U10618 ( .A(register__n6902), .Y(register__n6901) );
  BUFx2_ASAP7_75t_R register___U10619 ( .A(Reg_data[498]), .Y(register__n6902) );
  BUFx3_ASAP7_75t_R register___U10620 ( .A(register__net110087), .Y(register__net110086) );
  BUFx2_ASAP7_75t_R register___U10621 ( .A(Reg_data[491]), .Y(register__net110087) );
  BUFx4f_ASAP7_75t_R register___U10622 ( .A(register__net93753), .Y(register__net110088) );
  BUFx2_ASAP7_75t_R register___U10623 ( .A(register__net93753), .Y(register__net110090) );
  BUFx3_ASAP7_75t_R register___U10624 ( .A(register__net110083), .Y(register__net110082) );
  BUFx2_ASAP7_75t_R register___U10625 ( .A(Reg_data[486]), .Y(register__net110083) );
  BUFx3_ASAP7_75t_R register___U10626 ( .A(register__net110079), .Y(register__net110078) );
  BUFx2_ASAP7_75t_R register___U10627 ( .A(Reg_data[485]), .Y(register__net110079) );
  BUFx3_ASAP7_75t_R register___U10628 ( .A(register__n6904), .Y(register__n6903) );
  BUFx2_ASAP7_75t_R register___U10629 ( .A(Reg_data[484]), .Y(register__n6904) );
  BUFx3_ASAP7_75t_R register___U10630 ( .A(register__n6906), .Y(register__n6905) );
  BUFx2_ASAP7_75t_R register___U10631 ( .A(Reg_data[482]), .Y(register__n6906) );
  BUFx3_ASAP7_75t_R register___U10632 ( .A(register__n6908), .Y(register__n6907) );
  BUFx2_ASAP7_75t_R register___U10633 ( .A(Reg_data[480]), .Y(register__n6908) );
  BUFx4f_ASAP7_75t_R register___U10634 ( .A(register__n9294), .Y(register__n6909) );
  BUFx2_ASAP7_75t_R register___U10635 ( .A(register__n9294), .Y(register__n6910) );
  BUFx2_ASAP7_75t_R register___U10636 ( .A(register__n9294), .Y(register__n6911) );
  BUFx3_ASAP7_75t_R register___U10637 ( .A(register__n6913), .Y(register__n6912) );
  BUFx2_ASAP7_75t_R register___U10638 ( .A(Reg_data[501]), .Y(register__n6913) );
  BUFx4f_ASAP7_75t_R register___U10639 ( .A(register__n9386), .Y(register__n6914) );
  BUFx2_ASAP7_75t_R register___U10640 ( .A(register__n9386), .Y(register__n6915) );
  BUFx2_ASAP7_75t_R register___U10641 ( .A(register__n9386), .Y(register__n6916) );
  BUFx3_ASAP7_75t_R register___U10642 ( .A(register__n6918), .Y(register__n6917) );
  BUFx2_ASAP7_75t_R register___U10643 ( .A(Reg_data[617]), .Y(register__n6918) );
  BUFx3_ASAP7_75t_R register___U10644 ( .A(register__n6920), .Y(register__n6919) );
  BUFx2_ASAP7_75t_R register___U10645 ( .A(Reg_data[681]), .Y(register__n6920) );
  BUFx3_ASAP7_75t_R register___U10646 ( .A(register__n6922), .Y(register__n6921) );
  BUFx2_ASAP7_75t_R register___U10647 ( .A(Reg_data[415]), .Y(register__n6922) );
  BUFx4f_ASAP7_75t_R register___U10648 ( .A(register__n9776), .Y(register__n6923) );
  BUFx2_ASAP7_75t_R register___U10649 ( .A(register__n9776), .Y(register__n6924) );
  BUFx2_ASAP7_75t_R register___U10650 ( .A(register__n9776), .Y(register__n6925) );
  BUFx3_ASAP7_75t_R register___U10651 ( .A(register__net110029), .Y(register__net110028) );
  BUFx2_ASAP7_75t_R register___U10652 ( .A(Reg_data[376]), .Y(register__net110029) );
  BUFx3_ASAP7_75t_R register___U10653 ( .A(register__net110025), .Y(register__net110024) );
  BUFx2_ASAP7_75t_R register___U10654 ( .A(Reg_data[751]), .Y(register__net110025) );
  BUFx3_ASAP7_75t_R register___U10655 ( .A(register__net110021), .Y(register__net110020) );
  BUFx2_ASAP7_75t_R register___U10656 ( .A(Reg_data[79]), .Y(register__net110021) );
  BUFx3_ASAP7_75t_R register___U10657 ( .A(register__n6927), .Y(register__n6926) );
  BUFx2_ASAP7_75t_R register___U10658 ( .A(Reg_data[649]), .Y(register__n6927) );
  BUFx3_ASAP7_75t_R register___U10659 ( .A(register__n6929), .Y(register__n6928) );
  BUFx2_ASAP7_75t_R register___U10660 ( .A(Reg_data[670]), .Y(register__n6929) );
  BUFx3_ASAP7_75t_R register___U10661 ( .A(register__n10212), .Y(register__n6930) );
  BUFx4f_ASAP7_75t_R register___U10662 ( .A(register__n10212), .Y(register__n6931) );
  BUFx2_ASAP7_75t_R register___U10663 ( .A(register__n10212), .Y(register__n6932) );
  BUFx3_ASAP7_75t_R register___U10664 ( .A(register__n6934), .Y(register__n6933) );
  BUFx2_ASAP7_75t_R register___U10665 ( .A(Reg_data[654]), .Y(register__n6934) );
  BUFx3_ASAP7_75t_R register___U10666 ( .A(register__n6936), .Y(register__n6935) );
  BUFx2_ASAP7_75t_R register___U10667 ( .A(Reg_data[316]), .Y(register__n6936) );
  BUFx3_ASAP7_75t_R register___U10668 ( .A(register__n6938), .Y(register__n6937) );
  BUFx2_ASAP7_75t_R register___U10669 ( .A(Reg_data[940]), .Y(register__n6938) );
  BUFx3_ASAP7_75t_R register___U10670 ( .A(register__n6940), .Y(register__n6939) );
  BUFx2_ASAP7_75t_R register___U10671 ( .A(Reg_data[652]), .Y(register__n6940) );
  BUFx3_ASAP7_75t_R register___U10672 ( .A(register__n6942), .Y(register__n6941) );
  BUFx2_ASAP7_75t_R register___U10673 ( .A(Reg_data[915]), .Y(register__n6942) );
  BUFx2_ASAP7_75t_R register___U10674 ( .A(register__n9826), .Y(register__n6943) );
  BUFx2_ASAP7_75t_R register___U10675 ( .A(register__n9826), .Y(register__n6944) );
  BUFx4f_ASAP7_75t_R register___U10676 ( .A(register__n9826), .Y(register__n6945) );
  BUFx3_ASAP7_75t_R register___U10677 ( .A(register__n6947), .Y(register__n6946) );
  BUFx2_ASAP7_75t_R register___U10678 ( .A(Reg_data[723]), .Y(register__n6947) );
  BUFx3_ASAP7_75t_R register___U10679 ( .A(register__n10249), .Y(register__n6948) );
  BUFx2_ASAP7_75t_R register___U10680 ( .A(register__n10249), .Y(register__n6949) );
  BUFx4f_ASAP7_75t_R register___U10681 ( .A(register__n10249), .Y(register__n6950) );
  BUFx3_ASAP7_75t_R register___U10682 ( .A(register__n6952), .Y(register__n6951) );
  BUFx2_ASAP7_75t_R register___U10683 ( .A(Reg_data[851]), .Y(register__n6952) );
  BUFx3_ASAP7_75t_R register___U10684 ( .A(register__n6954), .Y(register__n6953) );
  BUFx2_ASAP7_75t_R register___U10685 ( .A(Reg_data[499]), .Y(register__n6954) );
  BUFx4f_ASAP7_75t_R register___U10686 ( .A(register__n9305), .Y(register__n6955) );
  BUFx2_ASAP7_75t_R register___U10687 ( .A(register__n9305), .Y(register__n6956) );
  BUFx2_ASAP7_75t_R register___U10688 ( .A(register__n9305), .Y(register__n6957) );
  BUFx3_ASAP7_75t_R register___U10689 ( .A(register__n6959), .Y(register__n6958) );
  BUFx2_ASAP7_75t_R register___U10690 ( .A(Reg_data[905]), .Y(register__n6959) );
  BUFx2_ASAP7_75t_R register___U10691 ( .A(register__n7682), .Y(register__n6960) );
  BUFx6f_ASAP7_75t_R register___U10692 ( .A(register__n7682), .Y(register__n6961) );
  BUFx3_ASAP7_75t_R register___U10693 ( .A(register__n6963), .Y(register__n6962) );
  BUFx2_ASAP7_75t_R register___U10694 ( .A(Reg_data[506]), .Y(register__n6963) );
  BUFx3_ASAP7_75t_R register___U10695 ( .A(register__n9311), .Y(register__n6964) );
  BUFx2_ASAP7_75t_R register___U10696 ( .A(register__n9311), .Y(register__n6965) );
  BUFx3_ASAP7_75t_R register___U10697 ( .A(register__n6968), .Y(register__n6967) );
  BUFx2_ASAP7_75t_R register___U10698 ( .A(Reg_data[241]), .Y(register__n6968) );
  BUFx3_ASAP7_75t_R register___U10699 ( .A(register__net109925), .Y(register__net109924) );
  BUFx2_ASAP7_75t_R register___U10700 ( .A(Reg_data[760]), .Y(register__net109925) );
  BUFx4f_ASAP7_75t_R register___U10701 ( .A(register__net90265), .Y(register__net109926) );
  BUFx2_ASAP7_75t_R register___U10702 ( .A(register__net90265), .Y(register__net109927) );
  BUFx3_ASAP7_75t_R register___U10703 ( .A(register__n6970), .Y(register__n6969) );
  BUFx2_ASAP7_75t_R register___U10704 ( .A(Reg_data[123]), .Y(register__n6970) );
  BUFx3_ASAP7_75t_R register___U10705 ( .A(register__n6972), .Y(register__n6971) );
  BUFx2_ASAP7_75t_R register___U10706 ( .A(Reg_data[379]), .Y(register__n6972) );
  BUFx4f_ASAP7_75t_R register___U10707 ( .A(register__n10507), .Y(register__n6973) );
  BUFx2_ASAP7_75t_R register___U10708 ( .A(register__n10507), .Y(register__n6974) );
  BUFx2_ASAP7_75t_R register___U10709 ( .A(register__n10507), .Y(register__n6975) );
  BUFx3_ASAP7_75t_R register___U10710 ( .A(register__net109907), .Y(register__net109906) );
  BUFx2_ASAP7_75t_R register___U10711 ( .A(Reg_data[381]), .Y(register__net109907) );
  BUFx3_ASAP7_75t_R register___U10712 ( .A(register__net109903), .Y(register__net109902) );
  BUFx2_ASAP7_75t_R register___U10713 ( .A(Reg_data[413]), .Y(register__net109903) );
  BUFx3_ASAP7_75t_R register___U10714 ( .A(register__net109899), .Y(register__net109898) );
  BUFx2_ASAP7_75t_R register___U10715 ( .A(Reg_data[445]), .Y(register__net109899) );
  BUFx3_ASAP7_75t_R register___U10716 ( .A(register__n6977), .Y(register__n6976) );
  BUFx2_ASAP7_75t_R register___U10717 ( .A(Reg_data[446]), .Y(register__n6977) );
  BUFx3_ASAP7_75t_R register___U10718 ( .A(register__n6979), .Y(register__n6978) );
  BUFx2_ASAP7_75t_R register___U10719 ( .A(Reg_data[494]), .Y(register__n6979) );
  BUFx2_ASAP7_75t_R register___U10720 ( .A(register__n9317), .Y(register__n6980) );
  BUFx2_ASAP7_75t_R register___U10721 ( .A(register__n9317), .Y(register__n6981) );
  BUFx4f_ASAP7_75t_R register___U10722 ( .A(register__n9317), .Y(register__n6982) );
  INVx2_ASAP7_75t_R register___U10723 ( .A(register__net97213), .Y(register__net109880) );
  BUFx6f_ASAP7_75t_R register___U10724 ( .A(register__net97214), .Y(register__net97213) );
  INVx2_ASAP7_75t_R register___U10725 ( .A(register__n8330), .Y(register__n11182) );
  BUFx6f_ASAP7_75t_R register___U10726 ( .A(register__n8331), .Y(register__n8330) );
  INVx2_ASAP7_75t_R register___U10727 ( .A(register__net94160), .Y(register__C6422_net59756) );
  BUFx6f_ASAP7_75t_R register___U10728 ( .A(register__net94161), .Y(register__net94160) );
  BUFx12f_ASAP7_75t_R register___U10729 ( .A(register__n12448), .Y(register__n12446) );
  BUFx4f_ASAP7_75t_R register___U10730 ( .A(register__n10662), .Y(register__n6984) );
  INVx2_ASAP7_75t_R register___U10731 ( .A(register__n8720), .Y(register__n10662) );
  BUFx6f_ASAP7_75t_R register___U10732 ( .A(register__n8721), .Y(register__n8720) );
  BUFx4f_ASAP7_75t_R register___U10733 ( .A(register__n10619), .Y(register__n6985) );
  INVx2_ASAP7_75t_R register___U10734 ( .A(register__n9209), .Y(register__n10619) );
  BUFx6f_ASAP7_75t_R register___U10735 ( .A(register__n9210), .Y(register__n9209) );
  INVx2_ASAP7_75t_R register___U10736 ( .A(register__net97193), .Y(register__net109852) );
  BUFx6f_ASAP7_75t_R register___U10737 ( .A(register__net97194), .Y(register__net97193) );
  OA22x2_ASAP7_75t_R register___U10738 ( .A1(register__n12021), .A2(register__n999), .B1(register__n10093), .B2(register__n972), 
        .Y(register__n13205) );
  INVx1_ASAP7_75t_R register___U10739 ( .A(register__n5970), .Y(register__n6986) );
  OA22x2_ASAP7_75t_R register___U10740 ( .A1(register__net63180), .A2(register__n7327), .B1(register__net88472), .B2(
        n11830), .Y(register__n12558) );
  INVx1_ASAP7_75t_R register___U10741 ( .A(register__n12558), .Y(register__n6989) );
  OA22x2_ASAP7_75t_R register___U10742 ( .A1(register__n12365), .A2(register__n1989), .B1(register__n10072), .B2(register__n3191), 
        .Y(register__n13341) );
  OA22x2_ASAP7_75t_R register___U10743 ( .A1(register__net64684), .A2(register__n2220), .B1(register__n10187), .B2(
        n11890), .Y(register__n12793) );
  INVx1_ASAP7_75t_R register___U10744 ( .A(register__n6248), .Y(register__n6990) );
  OA22x2_ASAP7_75t_R register___U10745 ( .A1(register__net64416), .A2(register__n1733), .B1(register__net89285), .B2(
        n3418), .Y(register__n13254) );
  OA22x2_ASAP7_75t_R register___U10746 ( .A1(register__net63324), .A2(register__n1706), .B1(register__n10253), .B2(
        n1739), .Y(register__n13246) );
  OA22x2_ASAP7_75t_R register___U10747 ( .A1(register__n12403), .A2(register__n1098), .B1(register__n10289), .B2(register__n535), 
        .Y(register__n12781) );
  OA22x2_ASAP7_75t_R register___U10748 ( .A1(register__n12394), .A2(register__n1988), .B1(register__n10301), .B2(register__n2155), 
        .Y(register__n13338) );
  OA22x2_ASAP7_75t_R register___U10749 ( .A1(register__net62834), .A2(register__n109), .B1(register__net89010), .B2(
        n11888), .Y(register__n12833) );
  INVx1_ASAP7_75t_R register___U10750 ( .A(register__n5097), .Y(register__n6992) );
  OA22x2_ASAP7_75t_R register___U10751 ( .A1(register__n12055), .A2(register__n1922), .B1(register__n7127), .B2(register__n1196), 
        .Y(register__n13107) );
  OA22x2_ASAP7_75t_R register___U10752 ( .A1(register__n11924), .A2(register__n982), .B1(register__n7479), .B2(register__n970), 
        .Y(register__n13207) );
  INVx1_ASAP7_75t_R register___U10753 ( .A(register__n13207), .Y(register__n6993) );
  OA22x2_ASAP7_75t_R register___U10754 ( .A1(register__net64016), .A2(register__n178), .B1(register__net103560), .B2(
        n206), .Y(register__n12677) );
  OA22x2_ASAP7_75t_R register___U10755 ( .A1(register__n12291), .A2(register__n187), .B1(register__n8162), .B2(register__n211), 
        .Y(register__n12673) );
  INVx1_ASAP7_75t_R register___U10756 ( .A(register__n4419), .Y(register__n6995) );
  OA22x2_ASAP7_75t_R register___U10757 ( .A1(register__n12082), .A2(register__n994), .B1(register__n7231), .B2(register__n973), 
        .Y(register__n13199) );
  OA22x2_ASAP7_75t_R register___U10758 ( .A1(register__n12229), .A2(register__n1922), .B1(register__n7147), .B2(register__n1212), 
        .Y(register__n13098) );
  INVx1_ASAP7_75t_R register___U10759 ( .A(register__net135334), .Y(register__net109782) );
  OA22x2_ASAP7_75t_R register___U10760 ( .A1(register__net64328), .A2(register__n1989), .B1(register__net89657), .B2(
        n5182), .Y(register__n13351) );
  OA22x2_ASAP7_75t_R register___U10761 ( .A1(register__net64664), .A2(register__n1988), .B1(register__n10160), .B2(
        n4953), .Y(register__n13354) );
  INVx2_ASAP7_75t_R register___U10762 ( .A(register__net62694), .Y(register__net62662) );
  OA22x2_ASAP7_75t_R register___U10763 ( .A1(register__n12454), .A2(register__n1006), .B1(register__n10195), .B2(register__n971), 
        .Y(register__n13178) );
  INVx1_ASAP7_75t_R register___U10764 ( .A(register__n10775), .Y(register__n7000) );
  INVx1_ASAP7_75t_R register___U10765 ( .A(register__n10777), .Y(register__n7002) );
  INVx1_ASAP7_75t_R register___U10766 ( .A(register__n5104), .Y(register__n7003) );
  INVx1_ASAP7_75t_R register___U10767 ( .A(register__n5106), .Y(register__n7004) );
  INVx1_ASAP7_75t_R register___U10768 ( .A(register__n5390), .Y(register__n7006) );
  INVx1_ASAP7_75t_R register___U10769 ( .A(register__n5736), .Y(register__n7007) );
  INVx1_ASAP7_75t_R register___U10770 ( .A(register__n4235), .Y(register__n7008) );
  INVx1_ASAP7_75t_R register___U10771 ( .A(register__n4237), .Y(register__n7009) );
  INVx1_ASAP7_75t_R register___U10772 ( .A(register__n4240), .Y(register__n7010) );
  INVx1_ASAP7_75t_R register___U10773 ( .A(register__n3091), .Y(register__n7011) );
  INVx1_ASAP7_75t_R register___U10774 ( .A(register__n3095), .Y(register__n7013) );
  INVx1_ASAP7_75t_R register___U10775 ( .A(register__n4348), .Y(register__n7014) );
  INVx1_ASAP7_75t_R register___U10776 ( .A(register__n4350), .Y(register__n7015) );
  AND4x1_ASAP7_75t_R register___U10777 ( .A(register__n1465), .B(register__n7014), .C(register__n7641), .D(register__n4352), .Y(
        n11449) );
  INVx1_ASAP7_75t_R register___U10778 ( .A(register__n5023), .Y(register__n7017) );
  INVx1_ASAP7_75t_R register___U10779 ( .A(register__n5025), .Y(register__n7018) );
  OA22x2_ASAP7_75t_R register___U10780 ( .A1(register__net64688), .A2(register__n175), .B1(register__n9720), .B2(register__n211), 
        .Y(register__n12685) );
  OA22x2_ASAP7_75t_R register___U10781 ( .A1(register__n12464), .A2(register__n7327), .B1(register__n9804), .B2(register__n3707), 
        .Y(register__n12554) );
  OA22x2_ASAP7_75t_R register___U10782 ( .A1(register__n12201), .A2(register__n2220), .B1(register__n9323), .B2(register__n7656), 
        .Y(register__n12786) );
  OA22x2_ASAP7_75t_R register___U10783 ( .A1(register__n12152), .A2(register__n116), .B1(register__n7376), .B2(register__n1658), 
        .Y(register__n12650) );
  OA22x2_ASAP7_75t_R register___U10784 ( .A1(register__n12205), .A2(register__n7327), .B1(register__n9585), .B2(register__n3539), 
        .Y(register__n12563) );
  OA22x2_ASAP7_75t_R register___U10785 ( .A1(register__net64860), .A2(register__n7327), .B1(register__net91069), .B2(
        n11832), .Y(register__n12573) );
  OA22x2_ASAP7_75t_R register___U10786 ( .A1(register__n11997), .A2(register__n7327), .B1(register__n5643), .B2(register__n4817), 
        .Y(register__n12576) );
  INVx1_ASAP7_75t_R register___U10787 ( .A(register__n5960), .Y(register__n7027) );
  OA22x2_ASAP7_75t_R register___U10788 ( .A1(register__n11934), .A2(register__n7327), .B1(register__n9595), .B2(register__n11833), 
        .Y(register__n12578) );
  OA22x2_ASAP7_75t_R register___U10789 ( .A1(register__n11933), .A2(register__n2119), .B1(register__n8706), .B2(register__n1682), 
        .Y(register__n12660) );
  INVx1_ASAP7_75t_R register___U10790 ( .A(register__n12660), .Y(register__n7029) );
  OA22x2_ASAP7_75t_R register___U10791 ( .A1(register__n11961), .A2(register__n181), .B1(register__n10485), .B2(register__n207), 
        .Y(register__n12690) );
  OA22x2_ASAP7_75t_R register___U10792 ( .A1(register__n12345), .A2(register__n109), .B1(register__n9955), .B2(register__n3021), 
        .Y(register__n12840) );
  INVx1_ASAP7_75t_R register___U10793 ( .A(register__n4868), .Y(register__n7030) );
  OA22x2_ASAP7_75t_R register___U10794 ( .A1(register__n11985), .A2(register__n1722), .B1(register__n6040), .B2(register__n1737), 
        .Y(register__n13261) );
  OA22x2_ASAP7_75t_R register___U10795 ( .A1(register__net63158), .A2(register__n1005), .B1(register__net93420), .B2(
        n975), .Y(register__n13183) );
  OA22x2_ASAP7_75t_R register___U10796 ( .A1(register__n12339), .A2(register__n998), .B1(register__n10511), .B2(register__n974), 
        .Y(register__n13187) );
  INVx1_ASAP7_75t_R register___U10797 ( .A(register__n5767), .Y(register__n7034) );
  INVx1_ASAP7_75t_R register___U10798 ( .A(register__n4401), .Y(register__n7035) );
  INVx1_ASAP7_75t_R register___U10799 ( .A(register__n4066), .Y(register__n7036) );
  OA22x2_ASAP7_75t_R register___U10800 ( .A1(register__n12153), .A2(register__n182), .B1(register__n9262), .B2(register__n219), 
        .Y(register__n12679) );
  INVx1_ASAP7_75t_R register___U10801 ( .A(register__n12679), .Y(register__n7037) );
  OA22x2_ASAP7_75t_R register___U10802 ( .A1(register__net64344), .A2(register__n702), .B1(register__net91367), .B2(
        n683), .Y(register__n13324) );
  OA22x2_ASAP7_75t_R register___U10803 ( .A1(register__net64336), .A2(register__n120), .B1(register__net97181), .B2(
        n1192), .Y(register__n13104) );
  OA22x2_ASAP7_75t_R register___U10804 ( .A1(register__net63008), .A2(register__n193), .B1(register__n8809), .B2(register__n206), 
        .Y(register__n12665) );
  INVx1_ASAP7_75t_R register___U10805 ( .A(register__n4407), .Y(register__n7039) );
  OA22x2_ASAP7_75t_R register___U10806 ( .A1(register__n3445), .A2(register__n1989), .B1(register__n10118), .B2(register__n11849), 
        .Y(register__n13348) );
  OA22x2_ASAP7_75t_R register___U10807 ( .A1(register__net129768), .A2(register__n1568), .B1(register__n9519), .B2(
        n1200), .Y(register__n13108) );
  INVx1_ASAP7_75t_R register___U10808 ( .A(register__n4072), .Y(register__n7040) );
  OA22x2_ASAP7_75t_R register___U10809 ( .A1(register__net64002), .A2(register__n1568), .B1(register__net93576), .B2(
        n1208), .Y(register__n13100) );
  INVx1_ASAP7_75t_R register___U10810 ( .A(register__n4074), .Y(register__n7041) );
  INVx1_ASAP7_75t_R register___U10811 ( .A(register__n5777), .Y(register__n7042) );
  OA22x2_ASAP7_75t_R register___U10812 ( .A1(register__n3186), .A2(register__n1922), .B1(register__n9559), .B2(register__n804), 
        .Y(register__n13089) );
  INVx1_ASAP7_75t_R register___U10813 ( .A(register__n5974), .Y(register__n7044) );
  OA22x2_ASAP7_75t_R register___U10814 ( .A1(register__net62828), .A2(register__n699), .B1(register__net91203), .B2(
        n675), .Y(register__n13308) );
  OA22x2_ASAP7_75t_R register___U10815 ( .A1(register__net64438), .A2(register__n105), .B1(register__net102363), .B2(
        n1661), .Y(register__n12653) );
  INVx1_ASAP7_75t_R register___U10816 ( .A(register__n5092), .Y(register__n7045) );
  OA22x2_ASAP7_75t_R register___U10817 ( .A1(register__n12293), .A2(register__n11915), .B1(register__register__n9828), .B2(register__n98), 
        .Y(register__n12562) );
  OA22x2_ASAP7_75t_R register___U10818 ( .A1(register__net63002), .A2(register__n109), .B1(register__n8821), .B2(register__n11801), .Y(register__n12835) );
  OA22x2_ASAP7_75t_R register___U10819 ( .A1(register__n12115), .A2(register__n118), .B1(register__n8740), .B2(register__n1205), 
        .Y(register__n13103) );
  INVx1_ASAP7_75t_R register___U10820 ( .A(register__n5791), .Y(register__n7046) );
  INVx4_ASAP7_75t_R register___U10821 ( .A(register__net63046), .Y(register__net63010) );
  OA22x2_ASAP7_75t_R register___U10822 ( .A1(register__net62986), .A2(register__n701), .B1(register__n10413), .B2(register__n696), 
        .Y(register__n13310) );
  INVx1_ASAP7_75t_R register___U10823 ( .A(register__n4543), .Y(register__n7047) );
  OA22x2_ASAP7_75t_R register___U10824 ( .A1(register__n12176), .A2(register__n117), .B1(register__n8829), .B2(register__n1675), 
        .Y(register__n12649) );
  INVx1_ASAP7_75t_R register___U10825 ( .A(register__n5099), .Y(register__n7048) );
  OA22x2_ASAP7_75t_R register___U10826 ( .A1(register__n12177), .A2(register__n7327), .B1(register__n5211), .B2(register__n3603), 
        .Y(register__n12565) );
  OA22x2_ASAP7_75t_R register___U10827 ( .A1(register__net62830), .A2(register__n101), .B1(register__net107858), .B2(
        n1919), .Y(register__n12951) );
  INVx1_ASAP7_75t_R register___U10828 ( .A(register__n13307), .Y(register__n7051) );
  INVx1_ASAP7_75t_R register___U10829 ( .A(register__n11267), .Y(register__n7053) );
  INVx1_ASAP7_75t_R register___U10830 ( .A(register__n3980), .Y(register__n7054) );
  INVx1_ASAP7_75t_R register___U10831 ( .A(register__n3982), .Y(register__n7055) );
  INVx1_ASAP7_75t_R register___U10832 ( .A(register__n4167), .Y(register__n7056) );
  INVx1_ASAP7_75t_R register___U10833 ( .A(register__n4169), .Y(register__n7057) );
  INVx1_ASAP7_75t_R register___U10834 ( .A(register__n4439), .Y(register__n7062) );
  INVx1_ASAP7_75t_R register___U10835 ( .A(register__n4730), .Y(register__n7065) );
  INVx1_ASAP7_75t_R register___U10836 ( .A(register__n4732), .Y(register__n7066) );
  INVx1_ASAP7_75t_R register___U10837 ( .A(register__n4914), .Y(register__n7067) );
  INVx1_ASAP7_75t_R register___U10838 ( .A(register__n4916), .Y(register__n7068) );
  INVx1_ASAP7_75t_R register___U10839 ( .A(register__n10560), .Y(register__n7070) );
  INVx1_ASAP7_75t_R register___U10840 ( .A(register__n3495), .Y(register__n7071) );
  INVx1_ASAP7_75t_R register___U10841 ( .A(register__n10557), .Y(register__n7072) );
  INVx1_ASAP7_75t_R register___U10842 ( .A(register__n4741), .Y(register__n7073) );
  OA22x2_ASAP7_75t_R register___U10843 ( .A1(register__n12376), .A2(register__net66574), .B1(register__n9435), .B2(
        n1674), .Y(register__n12641) );
  OA22x2_ASAP7_75t_R register___U10844 ( .A1(register__n12062), .A2(register__n111), .B1(register__n9439), .B2(register__n1681), 
        .Y(register__n12655) );
  OA22x2_ASAP7_75t_R register___U10845 ( .A1(register__net64774), .A2(register__n114), .B1(register__net91527), .B2(
        n1677), .Y(register__n12656) );
  INVx1_ASAP7_75t_R register___U10846 ( .A(register__n12656), .Y(register__n7075) );
  OA22x2_ASAP7_75t_R register___U10847 ( .A1(register__n11996), .A2(register__n116), .B1(register__n9443), .B2(register__n1680), 
        .Y(register__n12658) );
  OA22x2_ASAP7_75t_R register___U10848 ( .A1(register__n3373), .A2(register__n1092), .B1(register__n9680), .B2(register__n3350), 
        .Y(register__n13087) );
  OA22x2_ASAP7_75t_R register___U10849 ( .A1(register__n1911), .A2(register__n1922), .B1(register__n8827), .B2(register__n1204), 
        .Y(register__n13097) );
  OA22x2_ASAP7_75t_R register___U10850 ( .A1(register__net64836), .A2(register__n118), .B1(register__net96610), .B2(
        n1209), .Y(register__n13110) );
  OA22x2_ASAP7_75t_R register___U10851 ( .A1(register__register__n11954), .A2(register__n120), .B1(register__n9375), .B2(register__n1195), 
        .Y(register__n13114) );
  OA22x2_ASAP7_75t_R register___U10852 ( .A1(register__n12337), .A2(register__n699), .B1(register__n9489), .B2(register__n681), 
        .Y(register__n13315) );
  INVx1_ASAP7_75t_R register___U10853 ( .A(register__n4505), .Y(register__n7080) );
  OA22x2_ASAP7_75t_R register___U10854 ( .A1(register__n12254), .A2(register__n698), .B1(register__n9493), .B2(register__n682), 
        .Y(register__n13318) );
  INVx1_ASAP7_75t_R register___U10855 ( .A(register__n4060), .Y(register__n7081) );
  OA22x2_ASAP7_75t_R register___U10856 ( .A1(register__n5684), .A2(register__n698), .B1(register__n9495), .B2(register__n691), 
        .Y(register__n13320) );
  OA22x2_ASAP7_75t_R register___U10857 ( .A1(register__net64750), .A2(register__n701), .B1(register__net91395), .B2(
        n697), .Y(register__n13329) );
  INVx1_ASAP7_75t_R register___U10858 ( .A(register__n4062), .Y(register__n7082) );
  OA22x2_ASAP7_75t_R register___U10859 ( .A1(register__net64834), .A2(register__n699), .B1(register__net88949), .B2(
        n674), .Y(register__n13330) );
  OA22x2_ASAP7_75t_R register___U10860 ( .A1(register__net64922), .A2(register__n702), .B1(register__n10349), .B2(register__n676), 
        .Y(register__n13331) );
  OA22x2_ASAP7_75t_R register___U10861 ( .A1(register__n3723), .A2(register__n699), .B1(register__n9499), .B2(register__n693), 
        .Y(register__n13333) );
  INVx1_ASAP7_75t_R register___U10862 ( .A(register__n4064), .Y(register__n7083) );
  OA22x2_ASAP7_75t_R register___U10863 ( .A1(register__n11988), .A2(register__n118), .B1(register__n10345), .B2(register__n1199), 
        .Y(register__n13113) );
  INVx1_ASAP7_75t_R register___U10864 ( .A(register__n4094), .Y(register__n7084) );
  OA22x2_ASAP7_75t_R register___U10865 ( .A1(register__net63178), .A2(register__n1653), .B1(register__net88977), .B2(
        n1667), .Y(register__n12639) );
  OA22x2_ASAP7_75t_R register___U10866 ( .A1(register__n11950), .A2(register__n699), .B1(register__n10351), .B2(register__n692), 
        .Y(register__n13334) );
  OA22x2_ASAP7_75t_R register___U10867 ( .A1(register__n12228), .A2(register__n1755), .B1(register__n8771), .B2(register__n3336), 
        .Y(register__n13130) );
  INVx1_ASAP7_75t_R register___U10868 ( .A(register__net113159), .Y(register__net109215) );
  BUFx2_ASAP7_75t_R register___U10869 ( .A(Reg_data[855]), .Y(register__net109216) );
  BUFx3_ASAP7_75t_R register___U10870 ( .A(register__net109216), .Y(register__C6423_net61090) );
  BUFx2_ASAP7_75t_R register___U10871 ( .A(register__n10766), .Y(register__n7089) );
  BUFx2_ASAP7_75t_R register___U10872 ( .A(register__n11043), .Y(register__n7090) );
  BUFx2_ASAP7_75t_R register___U10873 ( .A(register__n11480), .Y(register__n7091) );
  BUFx2_ASAP7_75t_R register___U10874 ( .A(register__C6423_net60645), .Y(register__net108801) );
  BUFx2_ASAP7_75t_R register___U10875 ( .A(register__n11226), .Y(register__n7092) );
  BUFx2_ASAP7_75t_R register___U10876 ( .A(register__n11435), .Y(register__n7093) );
  INVx2_ASAP7_75t_R register___U10877 ( .A(register__n9483), .Y(register__n10575) );
  BUFx2_ASAP7_75t_R register___U10878 ( .A(register__n10529), .Y(register__n7094) );
  BUFx2_ASAP7_75t_R register___U10879 ( .A(register__n10936), .Y(register__n7095) );
  BUFx2_ASAP7_75t_R register___U10880 ( .A(register__n10866), .Y(register__n7096) );
  INVx2_ASAP7_75t_R register___U10881 ( .A(register__n9469), .Y(register__n11203) );
  INVx2_ASAP7_75t_R register___U10882 ( .A(register__n9459), .Y(register__n11567) );
  BUFx2_ASAP7_75t_R register___U10883 ( .A(register__n11392), .Y(register__n7097) );
  BUFx2_ASAP7_75t_R register___U10884 ( .A(register__n10682), .Y(register__n7098) );
  BUFx2_ASAP7_75t_R register___U10885 ( .A(register__n11104), .Y(register__n7099) );
  BUFx2_ASAP7_75t_R register___U10886 ( .A(register__n11350), .Y(register__n7100) );
  BUFx2_ASAP7_75t_R register___U10887 ( .A(register__C6422_net59959), .Y(register__net108770) );
  BUFx2_ASAP7_75t_R register___U10888 ( .A(register__n10890), .Y(register__n7101) );
  BUFx2_ASAP7_75t_R register___U10889 ( .A(register__n10739), .Y(register__n7102) );
  BUFx2_ASAP7_75t_R register___U10890 ( .A(register__n11412), .Y(register__n7103) );
  BUFx2_ASAP7_75t_R register___U10891 ( .A(register__n11707), .Y(register__n7104) );
  INVx2_ASAP7_75t_R register___U10892 ( .A(register__n10395), .Y(register__n11062) );
  BUFx2_ASAP7_75t_R register___U10893 ( .A(register__C6423_net61114), .Y(register__net108759) );
  BUFx2_ASAP7_75t_R register___U10894 ( .A(register__n11501), .Y(register__n7105) );
  BUFx2_ASAP7_75t_R register___U10895 ( .A(register__n11059), .Y(register__n7106) );
  BUFx2_ASAP7_75t_R register___U10896 ( .A(register__n11624), .Y(register__n7107) );
  BUFx2_ASAP7_75t_R register___U10897 ( .A(register__n11019), .Y(register__n7108) );
  INVx2_ASAP7_75t_R register___U10898 ( .A(register__n10385), .Y(register__n11105) );
  BUFx2_ASAP7_75t_R register___U10899 ( .A(register__C6422_net60326), .Y(register__net108748) );
  BUFx2_ASAP7_75t_R register___U10900 ( .A(register__n11372), .Y(register__n7109) );
  BUFx3_ASAP7_75t_R register___U10901 ( .A(register__n7111), .Y(register__n7110) );
  BUFx2_ASAP7_75t_R register___U10902 ( .A(register__n10967), .Y(register__n7111) );
  BUFx3_ASAP7_75t_R register___U10903 ( .A(register__n7113), .Y(register__n7112) );
  BUFx2_ASAP7_75t_R register___U10904 ( .A(register__n10710), .Y(register__n7113) );
  BUFx3_ASAP7_75t_R register___U10905 ( .A(register__n7115), .Y(register__n7114) );
  BUFx2_ASAP7_75t_R register___U10906 ( .A(register__n11033), .Y(register__n7115) );
  BUFx2_ASAP7_75t_R register___U10907 ( .A(register__n7121), .Y(register__n7120) );
  BUFx2_ASAP7_75t_R register___U10908 ( .A(register__n12842), .Y(register__n7121) );
  BUFx2_ASAP7_75t_R register___U10909 ( .A(register__n7123), .Y(register__n7122) );
  BUFx3_ASAP7_75t_R register___U10910 ( .A(register__n7714), .Y(register__n7124) );
  BUFx4f_ASAP7_75t_R register___U10911 ( .A(register__n7124), .Y(register__n8707) );
  BUFx2_ASAP7_75t_R register___U10912 ( .A(Reg_data[328]), .Y(register__n7125) );
  BUFx4f_ASAP7_75t_R register___U10913 ( .A(register__n7128), .Y(register__n7126) );
  BUFx6f_ASAP7_75t_R register___U10914 ( .A(register__n8686), .Y(register__n7128) );
  BUFx6f_ASAP7_75t_R register___U10915 ( .A(register__n7126), .Y(register__n10665) );
  BUFx4f_ASAP7_75t_R register___U10916 ( .A(register__n8687), .Y(register__n8686) );
  BUFx3_ASAP7_75t_R register___U10917 ( .A(register__n7125), .Y(register__n8687) );
  BUFx3_ASAP7_75t_R register___U10918 ( .A(register__net106198), .Y(register__net108339) );
  BUFx12f_ASAP7_75t_R register___U10919 ( .A(register__n10161), .Y(register__n7129) );
  BUFx3_ASAP7_75t_R register___U10920 ( .A(register__net98423), .Y(register__net108335) );
  BUFx3_ASAP7_75t_R register___U10921 ( .A(register__net98408), .Y(register__net108333) );
  BUFx3_ASAP7_75t_R register___U10922 ( .A(register__n7715), .Y(register__n7130) );
  BUFx4f_ASAP7_75t_R register___U10923 ( .A(register__n7130), .Y(register__n8733) );
  BUFx2_ASAP7_75t_R register___U10924 ( .A(Reg_data[787]), .Y(register__n7131) );
  BUFx2_ASAP7_75t_R register___U10925 ( .A(register__n7659), .Y(register__n7132) );
  BUFx4f_ASAP7_75t_R register___U10926 ( .A(register__n7659), .Y(register__n7133) );
  BUFx6f_ASAP7_75t_R register___U10927 ( .A(register__n7133), .Y(register__n11500) );
  BUFx4f_ASAP7_75t_R register___U10928 ( .A(register__n7660), .Y(register__n7659) );
  BUFx3_ASAP7_75t_R register___U10929 ( .A(register__n7131), .Y(register__n7660) );
  BUFx3_ASAP7_75t_R register___U10930 ( .A(register__n7565), .Y(register__n7134) );
  BUFx3_ASAP7_75t_R register___U10931 ( .A(register__n7727), .Y(register__n7135) );
  BUFx4f_ASAP7_75t_R register___U10932 ( .A(register__n7135), .Y(register__n9218) );
  BUFx3_ASAP7_75t_R register___U10933 ( .A(register__net103891), .Y(register__net108313) );
  BUFx4f_ASAP7_75t_R register___U10934 ( .A(register__net108313), .Y(register__net94145) );
  BUFx3_ASAP7_75t_R register___U10935 ( .A(register__net108239), .Y(register__net108238) );
  BUFx2_ASAP7_75t_R register___U10936 ( .A(Reg_data[773]), .Y(register__net108239) );
  BUFx4f_ASAP7_75t_R register___U10937 ( .A(register__net108238), .Y(register__net99941) );
  BUFx3_ASAP7_75t_R register___U10938 ( .A(register__n7137), .Y(register__n7136) );
  BUFx2_ASAP7_75t_R register___U10939 ( .A(Reg_data[272]), .Y(register__n7137) );
  BUFx4f_ASAP7_75t_R register___U10940 ( .A(register__n7136), .Y(register__n8719) );
  BUFx2_ASAP7_75t_R register___U10941 ( .A(Reg_data[99]), .Y(register__n7138) );
  BUFx6f_ASAP7_75t_R register___U10942 ( .A(register__n10047), .Y(register__n10046) );
  BUFx4f_ASAP7_75t_R register___U10943 ( .A(register__n6810), .Y(register__n10047) );
  BUFx2_ASAP7_75t_R register___U10944 ( .A(Reg_data[625]), .Y(register__n7139) );
  BUFx4f_ASAP7_75t_R register___U10945 ( .A(register__n10100), .Y(register__n7140) );
  BUFx2_ASAP7_75t_R register___U10946 ( .A(register__n10100), .Y(register__n7141) );
  BUFx3_ASAP7_75t_R register___U10947 ( .A(register__n10100), .Y(register__n7142) );
  BUFx6f_ASAP7_75t_R register___U10948 ( .A(register__n10101), .Y(register__n10100) );
  BUFx4f_ASAP7_75t_R register___U10949 ( .A(register__n6275), .Y(register__n10101) );
  BUFx3_ASAP7_75t_R register___U10950 ( .A(register__net108215), .Y(register__net108214) );
  BUFx2_ASAP7_75t_R register___U10951 ( .A(Reg_data[842]), .Y(register__net108215) );
  BUFx4f_ASAP7_75t_R register___U10952 ( .A(register__net108214), .Y(register__net102364) );
  BUFx3_ASAP7_75t_R register___U10953 ( .A(register__n7144), .Y(register__n7143) );
  BUFx2_ASAP7_75t_R register___U10954 ( .A(Reg_data[332]), .Y(register__n7144) );
  BUFx4f_ASAP7_75t_R register___U10955 ( .A(register__n7143), .Y(register__n8741) );
  BUFx3_ASAP7_75t_R register___U10956 ( .A(register__n7146), .Y(register__n7145) );
  BUFx2_ASAP7_75t_R register___U10957 ( .A(Reg_data[337]), .Y(register__n7146) );
  BUFx4f_ASAP7_75t_R register___U10958 ( .A(register__n8332), .Y(register__n7147) );
  BUFx4f_ASAP7_75t_R register___U10959 ( .A(register__n8332), .Y(register__n7148) );
  BUFx4f_ASAP7_75t_R register___U10960 ( .A(register__n7145), .Y(register__n8333) );
  INVx1_ASAP7_75t_R register___U10961 ( .A(register__n5562), .Y(register__n7149) );
  INVx1_ASAP7_75t_R register___U10962 ( .A(register__n5399), .Y(register__n7150) );
  INVx3_ASAP7_75t_R register___U10963 ( .A(register__n11967), .Y(register__n11950) );
  BUFx6f_ASAP7_75t_R register___U10964 ( .A(register__n9405), .Y(register__n11967) );
  BUFx12f_ASAP7_75t_R register___U10965 ( .A(register__net117948), .Y(register__net66316) );
  BUFx3_ASAP7_75t_R register___U10966 ( .A(register__net108119), .Y(register__net108118) );
  BUFx2_ASAP7_75t_R register___U10967 ( .A(Reg_data[902]), .Y(register__net108119) );
  BUFx3_ASAP7_75t_R register___U10968 ( .A(register__net108115), .Y(register__net108114) );
  BUFx2_ASAP7_75t_R register___U10969 ( .A(Reg_data[901]), .Y(register__net108115) );
  BUFx2_ASAP7_75t_R register___U10970 ( .A(Reg_data[744]), .Y(register__n7152) );
  BUFx3_ASAP7_75t_R register___U10971 ( .A(register__net108104), .Y(register__net108103) );
  BUFx2_ASAP7_75t_R register___U10972 ( .A(Reg_data[729]), .Y(register__net108104) );
  BUFx3_ASAP7_75t_R register___U10973 ( .A(register__net108100), .Y(register__net108099) );
  BUFx2_ASAP7_75t_R register___U10974 ( .A(Reg_data[709]), .Y(register__net108100) );
  BUFx3_ASAP7_75t_R register___U10975 ( .A(register__n7154), .Y(register__n7153) );
  BUFx2_ASAP7_75t_R register___U10976 ( .A(Reg_data[704]), .Y(register__n7154) );
  BUFx3_ASAP7_75t_R register___U10977 ( .A(register__n7156), .Y(register__n7155) );
  BUFx2_ASAP7_75t_R register___U10978 ( .A(Reg_data[690]), .Y(register__n7156) );
  BUFx3_ASAP7_75t_R register___U10979 ( .A(register__n7158), .Y(register__n7157) );
  BUFx2_ASAP7_75t_R register___U10980 ( .A(Reg_data[688]), .Y(register__n7158) );
  BUFx3_ASAP7_75t_R register___U10981 ( .A(register__n7160), .Y(register__n7159) );
  BUFx2_ASAP7_75t_R register___U10982 ( .A(Reg_data[676]), .Y(register__n7160) );
  BUFx3_ASAP7_75t_R register___U10983 ( .A(register__n7162), .Y(register__n7161) );
  BUFx2_ASAP7_75t_R register___U10984 ( .A(Reg_data[660]), .Y(register__n7162) );
  BUFx3_ASAP7_75t_R register___U10985 ( .A(register__n7164), .Y(register__n7163) );
  BUFx2_ASAP7_75t_R register___U10986 ( .A(Reg_data[656]), .Y(register__n7164) );
  BUFx3_ASAP7_75t_R register___U10987 ( .A(register__net108072), .Y(register__net108071) );
  BUFx2_ASAP7_75t_R register___U10988 ( .A(Reg_data[473]), .Y(register__net108072) );
  BUFx3_ASAP7_75t_R register___U10989 ( .A(register__net108068), .Y(register__net108067) );
  BUFx2_ASAP7_75t_R register___U10990 ( .A(Reg_data[453]), .Y(register__net108068) );
  BUFx3_ASAP7_75t_R register___U10991 ( .A(register__n7166), .Y(register__n7165) );
  BUFx2_ASAP7_75t_R register___U10992 ( .A(Reg_data[451]), .Y(register__n7166) );
  BUFx3_ASAP7_75t_R register___U10993 ( .A(register__n7168), .Y(register__n7167) );
  BUFx2_ASAP7_75t_R register___U10994 ( .A(Reg_data[418]), .Y(register__n7168) );
  BUFx3_ASAP7_75t_R register___U10995 ( .A(register__n7170), .Y(register__n7169) );
  BUFx2_ASAP7_75t_R register___U10996 ( .A(Reg_data[417]), .Y(register__n7170) );
  BUFx3_ASAP7_75t_R register___U10997 ( .A(register__n7172), .Y(register__n7171) );
  BUFx2_ASAP7_75t_R register___U10998 ( .A(Reg_data[416]), .Y(register__n7172) );
  BUFx3_ASAP7_75t_R register___U10999 ( .A(register__n7174), .Y(register__n7173) );
  BUFx2_ASAP7_75t_R register___U11000 ( .A(Reg_data[405]), .Y(register__n7174) );
  BUFx3_ASAP7_75t_R register___U11001 ( .A(register__n7176), .Y(register__n7175) );
  BUFx2_ASAP7_75t_R register___U11002 ( .A(Reg_data[386]), .Y(register__n7176) );
  BUFx3_ASAP7_75t_R register___U11003 ( .A(register__n7178), .Y(register__n7177) );
  BUFx2_ASAP7_75t_R register___U11004 ( .A(Reg_data[356]), .Y(register__n7178) );
  BUFx3_ASAP7_75t_R register___U11005 ( .A(register__net108036), .Y(register__net108035) );
  BUFx2_ASAP7_75t_R register___U11006 ( .A(Reg_data[25]), .Y(register__net108036) );
  BUFx3_ASAP7_75t_R register___U11007 ( .A(register__n7180), .Y(register__n7179) );
  BUFx2_ASAP7_75t_R register___U11008 ( .A(Reg_data[22]), .Y(register__n7180) );
  BUFx3_ASAP7_75t_R register___U11009 ( .A(register__net108028), .Y(register__net108027) );
  BUFx2_ASAP7_75t_R register___U11010 ( .A(Reg_data[249]), .Y(register__net108028) );
  BUFx3_ASAP7_75t_R register___U11011 ( .A(register__n7182), .Y(register__n7181) );
  BUFx2_ASAP7_75t_R register___U11012 ( .A(Reg_data[40]), .Y(register__n7182) );
  BUFx3_ASAP7_75t_R register___U11013 ( .A(register__net108020), .Y(register__net108019) );
  BUFx2_ASAP7_75t_R register___U11014 ( .A(Reg_data[747]), .Y(register__net108020) );
  BUFx3_ASAP7_75t_R register___U11015 ( .A(register__net108011), .Y(register__net108010) );
  BUFx2_ASAP7_75t_R register___U11016 ( .A(Reg_data[715]), .Y(register__net108011) );
  BUFx12f_ASAP7_75t_R register___U11017 ( .A(register__net108013), .Y(register__net89593) );
  BUFx12f_ASAP7_75t_R register___U11018 ( .A(register__net89594), .Y(register__net108013) );
  BUFx3_ASAP7_75t_R register___U11019 ( .A(register__n7184), .Y(register__n7183) );
  BUFx2_ASAP7_75t_R register___U11020 ( .A(Reg_data[634]), .Y(register__n7184) );
  BUFx3_ASAP7_75t_R register___U11021 ( .A(register__n7186), .Y(register__n7185) );
  BUFx2_ASAP7_75t_R register___U11022 ( .A(Reg_data[749]), .Y(register__n7186) );
  BUFx3_ASAP7_75t_R register___U11023 ( .A(register__n7188), .Y(register__n7187) );
  BUFx2_ASAP7_75t_R register___U11024 ( .A(Reg_data[411]), .Y(register__n7188) );
  BUFx3_ASAP7_75t_R register___U11025 ( .A(register__n7190), .Y(register__n7189) );
  BUFx2_ASAP7_75t_R register___U11026 ( .A(Reg_data[809]), .Y(register__n7190) );
  BUFx3_ASAP7_75t_R register___U11027 ( .A(register__n9772), .Y(register__n7191) );
  BUFx2_ASAP7_75t_R register___U11028 ( .A(register__n9772), .Y(register__n7192) );
  BUFx4f_ASAP7_75t_R register___U11029 ( .A(register__n9772), .Y(register__n7193) );
  BUFx3_ASAP7_75t_R register___U11030 ( .A(register__net107985), .Y(register__net107984) );
  BUFx2_ASAP7_75t_R register___U11031 ( .A(Reg_data[24]), .Y(register__net107985) );
  BUFx4f_ASAP7_75t_R register___U11032 ( .A(register__n6528), .Y(register__n7194) );
  BUFx2_ASAP7_75t_R register___U11033 ( .A(Reg_data[743]), .Y(register__n7195) );
  BUFx12f_ASAP7_75t_R register___U11034 ( .A(register__n9779), .Y(register__n9778) );
  BUFx6f_ASAP7_75t_R register___U11035 ( .A(register__n7194), .Y(register__n9779) );
  BUFx3_ASAP7_75t_R register___U11036 ( .A(register__n7197), .Y(register__n7196) );
  BUFx2_ASAP7_75t_R register___U11037 ( .A(Reg_data[318]), .Y(register__n7197) );
  BUFx3_ASAP7_75t_R register___U11038 ( .A(register__net107971), .Y(register__net107970) );
  BUFx2_ASAP7_75t_R register___U11039 ( .A(Reg_data[650]), .Y(register__net107971) );
  BUFx3_ASAP7_75t_R register___U11040 ( .A(register__n7199), .Y(register__n7198) );
  BUFx2_ASAP7_75t_R register___U11041 ( .A(Reg_data[60]), .Y(register__n7199) );
  BUFx3_ASAP7_75t_R register___U11042 ( .A(register__n7201), .Y(register__n7200) );
  BUFx2_ASAP7_75t_R register___U11043 ( .A(Reg_data[812]), .Y(register__n7201) );
  BUFx3_ASAP7_75t_R register___U11044 ( .A(register__n7203), .Y(register__n7202) );
  BUFx2_ASAP7_75t_R register___U11045 ( .A(Reg_data[172]), .Y(register__n7203) );
  BUFx3_ASAP7_75t_R register___U11046 ( .A(register__n7205), .Y(register__n7204) );
  BUFx2_ASAP7_75t_R register___U11047 ( .A(Reg_data[243]), .Y(register__n7205) );
  BUFx3_ASAP7_75t_R register___U11048 ( .A(register__n7207), .Y(register__n7206) );
  BUFx2_ASAP7_75t_R register___U11049 ( .A(Reg_data[531]), .Y(register__n7207) );
  BUFx3_ASAP7_75t_R register___U11050 ( .A(register__net107941), .Y(register__net107940) );
  BUFx2_ASAP7_75t_R register___U11051 ( .A(Reg_data[234]), .Y(register__net107941) );
  BUFx2_ASAP7_75t_R register___U11052 ( .A(register__net93396), .Y(register__net107943) );
  BUFx4f_ASAP7_75t_R register___U11053 ( .A(register__net93396), .Y(register__net107944) );
  BUFx4f_ASAP7_75t_R register___U11054 ( .A(register__n6046), .Y(register__n7208) );
  BUFx2_ASAP7_75t_R register___U11055 ( .A(Reg_data[759]), .Y(register__n7209) );
  BUFx12f_ASAP7_75t_R register___U11056 ( .A(register__n9831), .Y(register__n7210) );
  BUFx6f_ASAP7_75t_R register___U11057 ( .A(register__n7208), .Y(register__n9831) );
  BUFx3_ASAP7_75t_R register___U11058 ( .A(register__n7212), .Y(register__n7211) );
  BUFx2_ASAP7_75t_R register___U11059 ( .A(Reg_data[919]), .Y(register__n7212) );
  BUFx3_ASAP7_75t_R register___U11060 ( .A(register__n7214), .Y(register__n7213) );
  BUFx2_ASAP7_75t_R register___U11061 ( .A(Reg_data[535]), .Y(register__n7214) );
  BUFx3_ASAP7_75t_R register___U11062 ( .A(register__n10255), .Y(register__n7215) );
  BUFx2_ASAP7_75t_R register___U11063 ( .A(register__n10255), .Y(register__n7216) );
  BUFx4f_ASAP7_75t_R register___U11064 ( .A(register__n10255), .Y(register__n7217) );
  BUFx3_ASAP7_75t_R register___U11065 ( .A(register__n7219), .Y(register__n7218) );
  BUFx2_ASAP7_75t_R register___U11066 ( .A(Reg_data[667]), .Y(register__n7219) );
  BUFx3_ASAP7_75t_R register___U11067 ( .A(register__n8823), .Y(register__n7220) );
  BUFx2_ASAP7_75t_R register___U11068 ( .A(register__n8823), .Y(register__n7221) );
  BUFx4f_ASAP7_75t_R register___U11069 ( .A(register__n8823), .Y(register__n7222) );
  BUFx3_ASAP7_75t_R register___U11070 ( .A(register__n7224), .Y(register__n7223) );
  BUFx2_ASAP7_75t_R register___U11071 ( .A(Reg_data[699]), .Y(register__n7224) );
  BUFx3_ASAP7_75t_R register___U11072 ( .A(register__n7226), .Y(register__n7225) );
  BUFx2_ASAP7_75t_R register___U11073 ( .A(Reg_data[23]), .Y(register__n7226) );
  BUFx3_ASAP7_75t_R register___U11074 ( .A(register__n7228), .Y(register__n7227) );
  BUFx2_ASAP7_75t_R register___U11075 ( .A(Reg_data[233]), .Y(register__n7228) );
  BUFx2_ASAP7_75t_R register___U11076 ( .A(register__n10277), .Y(register__n7229) );
  BUFx2_ASAP7_75t_R register___U11077 ( .A(register__n10277), .Y(register__n7230) );
  BUFx4f_ASAP7_75t_R register___U11078 ( .A(register__n10277), .Y(register__n7231) );
  BUFx3_ASAP7_75t_R register___U11079 ( .A(register__n7233), .Y(register__n7232) );
  BUFx2_ASAP7_75t_R register___U11080 ( .A(Reg_data[474]), .Y(register__n7233) );
  BUFx3_ASAP7_75t_R register___U11081 ( .A(register__n7235), .Y(register__n7234) );
  BUFx2_ASAP7_75t_R register___U11082 ( .A(Reg_data[26]), .Y(register__n7235) );
  BUFx3_ASAP7_75t_R register___U11083 ( .A(register__n7237), .Y(register__n7236) );
  BUFx2_ASAP7_75t_R register___U11084 ( .A(Reg_data[209]), .Y(register__n7237) );
  BUFx3_ASAP7_75t_R register___U11085 ( .A(register__net107875), .Y(register__net107874) );
  BUFx2_ASAP7_75t_R register___U11086 ( .A(Reg_data[920]), .Y(register__net107875) );
  BUFx3_ASAP7_75t_R register___U11087 ( .A(register__net107871), .Y(register__net107870) );
  BUFx2_ASAP7_75t_R register___U11088 ( .A(Reg_data[696]), .Y(register__net107871) );
  BUFx3_ASAP7_75t_R register___U11089 ( .A(register__net107867), .Y(register__net107866) );
  BUFx2_ASAP7_75t_R register___U11090 ( .A(Reg_data[728]), .Y(register__net107867) );
  BUFx3_ASAP7_75t_R register___U11091 ( .A(register__net107857), .Y(register__net107856) );
  BUFx2_ASAP7_75t_R register___U11092 ( .A(Reg_data[509]), .Y(register__net107857) );
  BUFx2_ASAP7_75t_R register___U11093 ( .A(register__net93673), .Y(register__net107858) );
  BUFx3_ASAP7_75t_R register___U11094 ( .A(register__net93673), .Y(register__net107859) );
  BUFx3_ASAP7_75t_R register___U11095 ( .A(register__net107853), .Y(register__net107852) );
  BUFx2_ASAP7_75t_R register___U11096 ( .A(Reg_data[829]), .Y(register__net107853) );
  BUFx3_ASAP7_75t_R register___U11097 ( .A(register__n7239), .Y(register__n7238) );
  BUFx2_ASAP7_75t_R register___U11098 ( .A(Reg_data[764]), .Y(register__n7239) );
  BUFx3_ASAP7_75t_R register___U11099 ( .A(register__n7241), .Y(register__n7240) );
  BUFx2_ASAP7_75t_R register___U11100 ( .A(Reg_data[510]), .Y(register__n7241) );
  INVx2_ASAP7_75t_R register___U11101 ( .A(register__net97181), .Y(register__net107836) );
  BUFx6f_ASAP7_75t_R register___U11102 ( .A(register__net97182), .Y(register__net97181) );
  INVx2_ASAP7_75t_R register___U11103 ( .A(register__n12238), .Y(register__n12225) );
  BUFx4f_ASAP7_75t_R register___U11104 ( .A(register__n11456), .Y(register__n7242) );
  INVx2_ASAP7_75t_R register___U11105 ( .A(register__n7661), .Y(register__n11456) );
  BUFx6f_ASAP7_75t_R register___U11106 ( .A(register__n7662), .Y(register__n7661) );
  INVx2_ASAP7_75t_R register___U11107 ( .A(register__net94168), .Y(register__net107815) );
  BUFx6f_ASAP7_75t_R register___U11108 ( .A(register__net94169), .Y(register__net94168) );
  BUFx4f_ASAP7_75t_R register___U11109 ( .A(register__n10620), .Y(register__n7243) );
  INVx2_ASAP7_75t_R register___U11110 ( .A(register__n8722), .Y(register__n10620) );
  BUFx6f_ASAP7_75t_R register___U11111 ( .A(register__n8723), .Y(register__n8722) );
  BUFx4f_ASAP7_75t_R register___U11112 ( .A(register__n10555), .Y(register__n7244) );
  INVx2_ASAP7_75t_R register___U11113 ( .A(register__n7986), .Y(register__n10555) );
  BUFx6f_ASAP7_75t_R register___U11114 ( .A(register__n7987), .Y(register__n7986) );
  INVx2_ASAP7_75t_R register___U11115 ( .A(register__n8726), .Y(register__n10640) );
  BUFx6f_ASAP7_75t_R register___U11116 ( .A(register__n8727), .Y(register__n8726) );
  BUFx4f_ASAP7_75t_R register___U11117 ( .A(register__n11585), .Y(register__n7246) );
  INVx2_ASAP7_75t_R register___U11118 ( .A(register__n9213), .Y(register__n11585) );
  BUFx6f_ASAP7_75t_R register___U11119 ( .A(register__n9214), .Y(register__n9213) );
  BUFx4f_ASAP7_75t_R register___U11120 ( .A(register__n11328), .Y(register__n7247) );
  INVx2_ASAP7_75t_R register___U11121 ( .A(register__n8710), .Y(register__n11328) );
  BUFx6f_ASAP7_75t_R register___U11122 ( .A(register__n8711), .Y(register__n8710) );
  INVx2_ASAP7_75t_R register___U11123 ( .A(register__net97225), .Y(register__net107791) );
  BUFx6f_ASAP7_75t_R register___U11124 ( .A(register__net97226), .Y(register__net97225) );
  OA22x2_ASAP7_75t_R register___U11125 ( .A1(register__n11922), .A2(register__n399), .B1(register__n10050), .B2(register__n5642), 
        .Y(register__n13306) );
  OA22x2_ASAP7_75t_R register___U11126 ( .A1(register__n11962), .A2(register__n11900), .B1(register__n10499), .B2(register__n4842), .Y(register__n12635) );
  OA22x2_ASAP7_75t_R register___U11127 ( .A1(register__net64354), .A2(register__n1729), .B1(register__net89589), .B2(
        n3419), .Y(register__n13253) );
  OA22x2_ASAP7_75t_R register___U11128 ( .A1(register__net63346), .A2(register__n4267), .B1(register__n9832), .B2(register__n3385), .Y(register__n12613) );
  INVx1_ASAP7_75t_R register___U11129 ( .A(register__n4533), .Y(register__n7248) );
  OA22x2_ASAP7_75t_R register___U11130 ( .A1(register__net63340), .A2(register__n1098), .B1(register__n10261), .B2(
        n5356), .Y(register__n12784) );
  OA22x2_ASAP7_75t_R register___U11131 ( .A1(register__n12405), .A2(register__n177), .B1(register__n9853), .B2(register__n212), 
        .Y(register__n12666) );
  OA22x2_ASAP7_75t_R register___U11132 ( .A1(register__net64774), .A2(register__n4267), .B1(register__net95453), .B2(
        n3282), .Y(register__n12630) );
  INVx1_ASAP7_75t_R register___U11133 ( .A(register__n12630), .Y(register__n7250) );
  OA22x2_ASAP7_75t_R register___U11134 ( .A1(register__net64354), .A2(register__n4267), .B1(register__net95245), .B2(
        n11822), .Y(register__n12625) );
  OA22x2_ASAP7_75t_R register___U11135 ( .A1(register__n12175), .A2(register__n11816), .B1(register__n7395), .B2(register__n1594), 
        .Y(register__n12704) );
  OA22x2_ASAP7_75t_R register___U11136 ( .A1(register__net63178), .A2(register__n3119), .B1(register__net89845), .B2(
        n5500), .Y(register__n13291) );
  INVx1_ASAP7_75t_R register___U11137 ( .A(register__n6240), .Y(register__n7251) );
  OA22x2_ASAP7_75t_R register___U11138 ( .A1(register__net63178), .A2(register__n11900), .B1(register__net90761), .B2(
        n4268), .Y(register__n12611) );
  OA22x2_ASAP7_75t_R register___U11139 ( .A1(register__net64858), .A2(register__n4267), .B1(register__net90729), .B2(
        n3328), .Y(register__n12631) );
  INVx1_ASAP7_75t_R register___U11140 ( .A(register__n4399), .Y(register__n7252) );
  OA22x2_ASAP7_75t_R register___U11141 ( .A1(register__net64352), .A2(register__n109), .B1(register__net89661), .B2(
        n2960), .Y(register__n12849) );
  INVx1_ASAP7_75t_R register___U11142 ( .A(register__n4875), .Y(register__n7253) );
  OA22x2_ASAP7_75t_R register___U11143 ( .A1(register__n12152), .A2(register__n4267), .B1(register__n9748), .B2(register__n11904), 
        .Y(register__n12623) );
  INVx1_ASAP7_75t_R register___U11144 ( .A(register__n4667), .Y(register__n7254) );
  OA22x2_ASAP7_75t_R register___U11145 ( .A1(register__net64682), .A2(register__n109), .B1(register__n10155), .B2(register__n3473), .Y(register__n12853) );
  OA22x2_ASAP7_75t_R register___U11146 ( .A1(register__n12235), .A2(register__n189), .B1(register__n9770), .B2(register__n218), 
        .Y(register__n12675) );
  OA22x2_ASAP7_75t_R register___U11147 ( .A1(register__n12453), .A2(register__n1716), .B1(register__n10203), .B2(register__n11753), .Y(register__n13240) );
  INVx1_ASAP7_75t_R register___U11148 ( .A(register__n6797), .Y(register__n7256) );
  OA22x2_ASAP7_75t_R register___U11149 ( .A1(register__n12460), .A2(register__n2220), .B1(register__n10216), .B2(register__n11804), .Y(register__n12777) );
  BUFx12f_ASAP7_75t_R register___U11150 ( .A(register__net112578), .Y(register__C6422_net69812) );
  BUFx6f_ASAP7_75t_R register___U11151 ( .A(register__n12448), .Y(register__n12445) );
  INVx1_ASAP7_75t_R register___U11152 ( .A(register__n3849), .Y(register__n7260) );
  INVx1_ASAP7_75t_R register___U11153 ( .A(register__n5395), .Y(register__n7261) );
  INVx1_ASAP7_75t_R register___U11154 ( .A(register__n4052), .Y(register__n7262) );
  AO22x1_ASAP7_75t_R register___U11155 ( .A1(register__n9299), .A2(register__C6423_net61318), .B1(register__n10199), 
        .B2(register__n1451), .Y(register__n11690) );
  INVx1_ASAP7_75t_R register___U11156 ( .A(register__n4288), .Y(register__n7263) );
  INVx1_ASAP7_75t_R register___U11157 ( .A(register__n4317), .Y(register__n7264) );
  INVx1_ASAP7_75t_R register___U11158 ( .A(register__n4320), .Y(register__n7265) );
  INVx1_ASAP7_75t_R register___U11159 ( .A(register__n4705), .Y(register__n7269) );
  OA22x2_ASAP7_75t_R register___U11160 ( .A1(register__n12311), .A2(register__n399), .B1(register__n10036), .B2(register__n3380), 
        .Y(register__n13296) );
  OA22x2_ASAP7_75t_R register___U11161 ( .A1(register__net64352), .A2(register__n183), .B1(register__net90713), .B2(
        n209), .Y(register__n12681) );
  INVx1_ASAP7_75t_R register___U11162 ( .A(register__n4300), .Y(register__n7277) );
  OA22x2_ASAP7_75t_R register___U11163 ( .A1(register__net129768), .A2(register__n3119), .B1(register__n10096), .B2(
        n3326), .Y(register__n13303) );
  INVx1_ASAP7_75t_R register___U11164 ( .A(register__n6500), .Y(register__n7278) );
  OA22x2_ASAP7_75t_R register___U11165 ( .A1(register__net64018), .A2(register__n4267), .B1(register__net90689), .B2(
        n3480), .Y(register__n12621) );
  INVx1_ASAP7_75t_R register___U11166 ( .A(register__n5574), .Y(register__n7279) );
  OA22x2_ASAP7_75t_R register___U11167 ( .A1(register__n12452), .A2(register__n399), .B1(register__n8376), .B2(register__n5343), 
        .Y(register__n13286) );
  INVx1_ASAP7_75t_R register___U11168 ( .A(register__n4879), .Y(register__n7280) );
  OA22x2_ASAP7_75t_R register___U11169 ( .A1(register__n12114), .A2(register__n4033), .B1(register__n9736), .B2(register__n7050), 
        .Y(register__n12540) );
  OA22x2_ASAP7_75t_R register___U11170 ( .A1(register__n4596), .A2(register__n4033), .B1(register__n9250), .B2(register__n3361), 
        .Y(register__n12532) );
  OA22x2_ASAP7_75t_R register___U11171 ( .A1(register__n12064), .A2(register__n4033), .B1(register__n10477), .B2(register__n3737), 
        .Y(register__n12544) );
  INVx1_ASAP7_75t_R register___U11172 ( .A(register__n3760), .Y(register__n7282) );
  OA22x2_ASAP7_75t_R register___U11173 ( .A1(register__n12029), .A2(register__n189), .B1(register__n210), .B2(register__n9615), 
        .Y(register__n12688) );
  OA22x2_ASAP7_75t_R register___U11174 ( .A1(register__net63172), .A2(register__n2220), .B1(register__net93440), .B2(
        n3306), .Y(register__n12782) );
  OA22x2_ASAP7_75t_R register___U11175 ( .A1(register__n12059), .A2(register__n1098), .B1(register__n9935), .B2(register__n11808), 
        .Y(register__n12792) );
  INVx4_ASAP7_75t_R register___U11176 ( .A(register__n12072), .Y(register__n12059) );
  OA22x2_ASAP7_75t_R register___U11177 ( .A1(register__n11930), .A2(register__n2220), .B1(register__n9941), .B2(register__n3413), 
        .Y(register__n12799) );
  OA22x2_ASAP7_75t_R register___U11178 ( .A1(register__net63178), .A2(register__n109), .B1(register__net90061), .B2(
        n3673), .Y(register__n12836) );
  OA22x2_ASAP7_75t_R register___U11179 ( .A1(register__n11929), .A2(register__n109), .B1(register__n9967), .B2(register__n1474), 
        .Y(register__n12858) );
  OA22x2_ASAP7_75t_R register___U11180 ( .A1(register__net64752), .A2(register__n1732), .B1(register__net112730), .B2(
        n11871), .Y(register__n13258) );
  OA22x2_ASAP7_75t_R register___U11181 ( .A1(register__net64836), .A2(register__n1704), .B1(register__net89909), .B2(
        n5170), .Y(register__n13259) );
  OA22x2_ASAP7_75t_R register___U11182 ( .A1(register__net64442), .A2(register__n4033), .B1(register__net93805), .B2(
        n11837), .Y(register__n12542) );
  OA22x2_ASAP7_75t_R register___U11183 ( .A1(register__net64012), .A2(register__n2220), .B1(register__net89641), .B2(
        n4632), .Y(register__n12787) );
  OA22x2_ASAP7_75t_R register___U11184 ( .A1(register__n12459), .A2(register__n109), .B1(register__n10104), .B2(register__n11886), 
        .Y(register__n12832) );
  OA22x2_ASAP7_75t_R register___U11185 ( .A1(register__n12404), .A2(register__n4033), .B1(register__n9347), .B2(register__n11918), 
        .Y(register__n12527) );
  INVx1_ASAP7_75t_R register___U11186 ( .A(register__n5972), .Y(register__n7289) );
  OA22x2_ASAP7_75t_R register___U11187 ( .A1(register__net63008), .A2(register__n4269), .B1(register__n9535), .B2(register__n1599), .Y(register__n12694) );
  OA22x2_ASAP7_75t_R register___U11188 ( .A1(register__net62986), .A2(register__n399), .B1(register__n10323), .B2(register__n5341), .Y(register__n13289) );
  INVx1_ASAP7_75t_R register___U11189 ( .A(register__n5981), .Y(register__n7290) );
  OA22x2_ASAP7_75t_R register___U11190 ( .A1(register__net62990), .A2(register__n1002), .B1(register__n8354), .B2(register__n972), 
        .Y(register__n13181) );
  OA22x2_ASAP7_75t_R register___U11191 ( .A1(register__n12375), .A2(register__n176), .B1(register__n6837), .B2(register__n221), 
        .Y(register__n12670) );
  INVx1_ASAP7_75t_R register___U11192 ( .A(register__n12670), .Y(register__n7291) );
  OA22x2_ASAP7_75t_R register___U11193 ( .A1(register__net63156), .A2(register__n1730), .B1(register__net119539), .B2(
        n1715), .Y(register__n13244) );
  INVx1_ASAP7_75t_R register___U11194 ( .A(register__n13244), .Y(register__n7292) );
  OA22x2_ASAP7_75t_R register___U11195 ( .A1(register__n12172), .A2(register__n109), .B1(register__n6876), .B2(register__n3674), 
        .Y(register__n12846) );
  INVx1_ASAP7_75t_R register___U11196 ( .A(register__n4877), .Y(register__n7293) );
  OA22x2_ASAP7_75t_R register___U11197 ( .A1(register__net62988), .A2(register__n1727), .B1(register__n10267), .B2(
        n1728), .Y(register__n13242) );
  OA22x2_ASAP7_75t_R register___U11198 ( .A1(register__n12462), .A2(register__n3022), .B1(register__n10387), .B2(register__n1587), 
        .Y(register__n12692) );
  INVx1_ASAP7_75t_R register___U11199 ( .A(register__n5785), .Y(register__n7294) );
  BUFx12f_ASAP7_75t_R register___U11200 ( .A(register__n12308), .Y(register__n7295) );
  BUFx12f_ASAP7_75t_R register___U11201 ( .A(register__n12308), .Y(register__n7296) );
  BUFx6f_ASAP7_75t_R register___U11202 ( .A(register__n3844), .Y(register__n12297) );
  BUFx6f_ASAP7_75t_R register___U11203 ( .A(register__n3446), .Y(register__n12298) );
  BUFx6f_ASAP7_75t_R register___U11204 ( .A(register__n3672), .Y(register__n12296) );
  BUFx12f_ASAP7_75t_R register___U11205 ( .A(register__n7295), .Y(register__n12294) );
  INVx1_ASAP7_75t_R register___U11206 ( .A(register__n4898), .Y(register__n7297) );
  INVx1_ASAP7_75t_R register___U11207 ( .A(register__n4901), .Y(register__n7298) );
  INVx1_ASAP7_75t_R register___U11208 ( .A(register__n4903), .Y(register__n7299) );
  INVx1_ASAP7_75t_R register___U11209 ( .A(register__n4694), .Y(register__n7301) );
  INVx1_ASAP7_75t_R register___U11210 ( .A(register__n4696), .Y(register__n7302) );
  AO22x2_ASAP7_75t_R register___U11211 ( .A1(register__n9254), .A2(register__net128122), .B1(register__n10058), .B2(
        n2000), .Y(register__n11248) );
  INVx1_ASAP7_75t_R register___U11212 ( .A(register__n4610), .Y(register__n7307) );
  INVx1_ASAP7_75t_R register___U11213 ( .A(register__n3099), .Y(register__n7309) );
  INVx1_ASAP7_75t_R register___U11214 ( .A(register__n3101), .Y(register__n7310) );
  INVx1_ASAP7_75t_R register___U11215 ( .A(register__n4342), .Y(register__n7311) );
  INVx1_ASAP7_75t_R register___U11216 ( .A(register__n4252), .Y(register__n7315) );
  INVx1_ASAP7_75t_R register___U11217 ( .A(register__n4254), .Y(register__n7316) );
  INVx1_ASAP7_75t_R register___U11218 ( .A(register__n2975), .Y(register__n7318) );
  INVx1_ASAP7_75t_R register___U11219 ( .A(register__n2978), .Y(register__n7319) );
  INVx1_ASAP7_75t_R register___U11220 ( .A(register__n2980), .Y(register__n7320) );
  OA22x2_ASAP7_75t_R register___U11221 ( .A1(register__n12260), .A2(register__n3022), .B1(register__n9449), .B2(register__n1603), 
        .Y(register__n12701) );
  OA22x2_ASAP7_75t_R register___U11222 ( .A1(register__net64772), .A2(register__n3022), .B1(register__net91495), .B2(
        n1591), .Y(register__n12711) );
  OA22x2_ASAP7_75t_R register___U11223 ( .A1(register__n11995), .A2(register__n11816), .B1(register__n9455), .B2(register__n1597), 
        .Y(register__n12715) );
  OA22x2_ASAP7_75t_R register___U11224 ( .A1(register__n1019), .A2(register__n1409), .B1(register__n9427), .B2(register__n11749), 
        .Y(register__n13282) );
  OA22x2_ASAP7_75t_R register___U11225 ( .A1(register__net132881), .A2(register__n4033), .B1(register__net93468), .B2(
        n11843), .Y(register__n12524) );
  INVx1_ASAP7_75t_R register___U11226 ( .A(register__n12524), .Y(register__n7325) );
  OA22x2_ASAP7_75t_R register___U11227 ( .A1(register__net64838), .A2(register__n101), .B1(register__net93737), .B2(
        n11773), .Y(register__n12974) );
  INVx1_ASAP7_75t_R register___U11228 ( .A(register__n2915), .Y(register__n7326) );
  OA22x2_ASAP7_75t_R register___U11229 ( .A1(register__n11961), .A2(register__n2935), .B1(register__n10339), .B2(register__n1604), 
        .Y(register__n12716) );
  BUFx4f_ASAP7_75t_R register___U11230 ( .A(register__net122349), .Y(register__net106940) );
  BUFx6f_ASAP7_75t_R register___U11231 ( .A(register__n7338), .Y(register__n7337) );
  BUFx4f_ASAP7_75t_R register___U11232 ( .A(register__n6092), .Y(register__n7338) );
  BUFx2_ASAP7_75t_R register___U11233 ( .A(register__C6423_net60643), .Y(register__net106698) );
  BUFx2_ASAP7_75t_R register___U11234 ( .A(register__n10597), .Y(register__n7339) );
  BUFx2_ASAP7_75t_R register___U11235 ( .A(register__n11567), .Y(register__n7340) );
  BUFx2_ASAP7_75t_R register___U11236 ( .A(register__n11225), .Y(register__n7341) );
  BUFx2_ASAP7_75t_R register___U11237 ( .A(register__n10957), .Y(register__n7342) );
  BUFx2_ASAP7_75t_R register___U11238 ( .A(register__n10763), .Y(register__n7343) );
  BUFx2_ASAP7_75t_R register___U11239 ( .A(register__n11393), .Y(register__n7344) );
  BUFx2_ASAP7_75t_R register___U11240 ( .A(register__n11105), .Y(register__n7345) );
  BUFx2_ASAP7_75t_R register___U11241 ( .A(register__n11644), .Y(register__n7346) );
  BUFx2_ASAP7_75t_R register___U11242 ( .A(register__n11041), .Y(register__n7347) );
  BUFx3_ASAP7_75t_R register___U11243 ( .A(register__n7349), .Y(register__n7348) );
  BUFx2_ASAP7_75t_R register___U11244 ( .A(register__n10988), .Y(register__n7349) );
  BUFx2_ASAP7_75t_R register___U11245 ( .A(register__n7357), .Y(register__n7356) );
  BUFx2_ASAP7_75t_R register___U11246 ( .A(register__n13117), .Y(register__n7357) );
  BUFx6f_ASAP7_75t_R register___U11247 ( .A(register__n7954), .Y(register__n10916) );
  BUFx3_ASAP7_75t_R register___U11248 ( .A(register__n10573), .Y(register__n7358) );
  BUFx3_ASAP7_75t_R register___U11249 ( .A(register__n7360), .Y(register__n7359) );
  BUFx3_ASAP7_75t_R register___U11250 ( .A(register__n10571), .Y(register__n7361) );
  BUFx4f_ASAP7_75t_R register___U11251 ( .A(register__n7361), .Y(register__n9189) );
  INVx2_ASAP7_75t_R register___U11252 ( .A(register__n9189), .Y(register__n7362) );
  BUFx3_ASAP7_75t_R register___U11253 ( .A(register__n7366), .Y(register__n7365) );
  BUFx2_ASAP7_75t_R register___U11254 ( .A(register__n11661), .Y(register__n7366) );
  BUFx3_ASAP7_75t_R register___U11255 ( .A(register__n7368), .Y(register__n7367) );
  BUFx2_ASAP7_75t_R register___U11256 ( .A(register__n11660), .Y(register__n7368) );
  BUFx4f_ASAP7_75t_R register___U11257 ( .A(register__n7367), .Y(register__n9238) );
  INVx2_ASAP7_75t_R register___U11258 ( .A(register__n9238), .Y(register__n7369) );
  BUFx12f_ASAP7_75t_R register___U11259 ( .A(register__n10009), .Y(register__n7370) );
  BUFx3_ASAP7_75t_R register___U11260 ( .A(register__n8028), .Y(register__n7371) );
  BUFx3_ASAP7_75t_R register___U11261 ( .A(register__n8032), .Y(register__n7372) );
  BUFx3_ASAP7_75t_R register___U11262 ( .A(register__net101448), .Y(register__net106320) );
  BUFx3_ASAP7_75t_R register___U11263 ( .A(register__n8034), .Y(register__n7373) );
  BUFx12f_ASAP7_75t_R register___U11264 ( .A(register__net89794), .Y(register__net89793) );
  BUFx3_ASAP7_75t_R register___U11265 ( .A(register__net101217), .Y(register__net106314) );
  BUFx3_ASAP7_75t_R register___U11266 ( .A(register__n8996), .Y(register__n7374) );
  BUFx3_ASAP7_75t_R register___U11267 ( .A(register__net103939), .Y(register__net106310) );
  BUFx2_ASAP7_75t_R register___U11268 ( .A(Reg_data[845]), .Y(register__n7375) );
  BUFx2_ASAP7_75t_R register___U11269 ( .A(register__n8282), .Y(register__n7376) );
  BUFx4f_ASAP7_75t_R register___U11270 ( .A(register__n8282), .Y(register__n7377) );
  BUFx6f_ASAP7_75t_R register___U11271 ( .A(register__n7377), .Y(register__n10765) );
  BUFx4f_ASAP7_75t_R register___U11272 ( .A(register__n8283), .Y(register__n8282) );
  BUFx3_ASAP7_75t_R register___U11273 ( .A(register__n7375), .Y(register__n8283) );
  BUFx12f_ASAP7_75t_R register___U11274 ( .A(register__n10204), .Y(register__n7378) );
  BUFx3_ASAP7_75t_R register___U11275 ( .A(register__net101056), .Y(register__net106297) );
  BUFx3_ASAP7_75t_R register___U11276 ( .A(register__net103924), .Y(register__net106295) );
  BUFx3_ASAP7_75t_R register___U11277 ( .A(register__net103440), .Y(register__net106293) );
  BUFx3_ASAP7_75t_R register___U11278 ( .A(register__n7722), .Y(register__n7379) );
  BUFx2_ASAP7_75t_R register___U11279 ( .A(Reg_data[836]), .Y(register__net106240) );
  BUFx3_ASAP7_75t_R register___U11280 ( .A(register__net106236), .Y(register__net106235) );
  BUFx2_ASAP7_75t_R register___U11281 ( .A(Reg_data[793]), .Y(register__net106236) );
  BUFx4f_ASAP7_75t_R register___U11282 ( .A(register__net106235), .Y(register__net94177) );
  BUFx3_ASAP7_75t_R register___U11283 ( .A(register__n7381), .Y(register__n7380) );
  BUFx2_ASAP7_75t_R register___U11284 ( .A(Reg_data[576]), .Y(register__n7381) );
  BUFx4f_ASAP7_75t_R register___U11285 ( .A(register__n7380), .Y(register__n8715) );
  BUFx2_ASAP7_75t_R register___U11286 ( .A(Reg_data[345]), .Y(register__net106228) );
  BUFx3_ASAP7_75t_R register___U11287 ( .A(register__n7383), .Y(register__n7382) );
  BUFx2_ASAP7_75t_R register___U11288 ( .A(Reg_data[341]), .Y(register__n7383) );
  BUFx4f_ASAP7_75t_R register___U11289 ( .A(register__n7382), .Y(register__n8717) );
  BUFx3_ASAP7_75t_R register___U11290 ( .A(register__n7385), .Y(register__n7384) );
  BUFx2_ASAP7_75t_R register___U11291 ( .A(Reg_data[276]), .Y(register__n7385) );
  BUFx4f_ASAP7_75t_R register___U11292 ( .A(register__n7384), .Y(register__n9212) );
  BUFx3_ASAP7_75t_R register___U11293 ( .A(register__net106214), .Y(register__net106213) );
  BUFx2_ASAP7_75t_R register___U11294 ( .A(Reg_data[262]), .Y(register__net106214) );
  BUFx4f_ASAP7_75t_R register___U11295 ( .A(register__net106213), .Y(register__net97198) );
  BUFx2_ASAP7_75t_R register___U11296 ( .A(Reg_data[260]), .Y(register__n7386) );
  BUFx2_ASAP7_75t_R register___U11297 ( .A(Reg_data[843]), .Y(register__net106198) );
  BUFx4f_ASAP7_75t_R register___U11298 ( .A(register__net106202), .Y(register__net106199) );
  BUFx6f_ASAP7_75t_R register___U11299 ( .A(register__net106201), .Y(register__net106200) );
  BUFx6f_ASAP7_75t_R register___U11300 ( .A(register__net102367), .Y(register__net106201) );
  BUFx3_ASAP7_75t_R register___U11301 ( .A(register__net102367), .Y(register__net106202) );
  BUFx6f_ASAP7_75t_R register___U11302 ( .A(register__net102368), .Y(register__net102367) );
  BUFx4f_ASAP7_75t_R register___U11303 ( .A(register__net108339), .Y(register__net102368) );
  BUFx3_ASAP7_75t_R register___U11304 ( .A(register__net106194), .Y(register__net106193) );
  BUFx2_ASAP7_75t_R register___U11305 ( .A(Reg_data[778]), .Y(register__net106194) );
  BUFx4f_ASAP7_75t_R register___U11306 ( .A(register__net106193), .Y(register__net97178) );
  BUFx2_ASAP7_75t_R register___U11307 ( .A(Reg_data[403]), .Y(register__n7387) );
  BUFx6f_ASAP7_75t_R register___U11308 ( .A(register__n9761), .Y(register__n9760) );
  BUFx4f_ASAP7_75t_R register___U11309 ( .A(register__n5511), .Y(register__n9761) );
  BUFx2_ASAP7_75t_R register___U11310 ( .A(Reg_data[263]), .Y(register__n7388) );
  BUFx2_ASAP7_75t_R register___U11311 ( .A(Reg_data[479]), .Y(register__n7389) );
  BUFx2_ASAP7_75t_R register___U11312 ( .A(register__n10438), .Y(register__n7390) );
  BUFx3_ASAP7_75t_R register___U11313 ( .A(register__n10438), .Y(register__n7391) );
  BUFx4f_ASAP7_75t_R register___U11314 ( .A(register__n10438), .Y(register__n7392) );
  BUFx6f_ASAP7_75t_R register___U11315 ( .A(register__n10439), .Y(register__n10438) );
  BUFx4f_ASAP7_75t_R register___U11316 ( .A(register__n5046), .Y(register__n10439) );
  BUFx3_ASAP7_75t_R register___U11317 ( .A(register__net106173), .Y(register__net106172) );
  BUFx2_ASAP7_75t_R register___U11318 ( .A(Reg_data[344]), .Y(register__net106173) );
  BUFx4f_ASAP7_75t_R register___U11319 ( .A(register__net106172), .Y(register__net97161) );
  BUFx3_ASAP7_75t_R register___U11320 ( .A(register__n7394), .Y(register__n7393) );
  BUFx2_ASAP7_75t_R register___U11321 ( .A(Reg_data[782]), .Y(register__n7394) );
  BUFx4f_ASAP7_75t_R register___U11322 ( .A(register__n8730), .Y(register__n7395) );
  BUFx4f_ASAP7_75t_R register___U11323 ( .A(register__n8730), .Y(register__n7396) );
  BUFx4f_ASAP7_75t_R register___U11324 ( .A(register__n7393), .Y(register__n8731) );
  BUFx3_ASAP7_75t_R register___U11325 ( .A(register__net106155), .Y(register__net106154) );
  BUFx2_ASAP7_75t_R register___U11326 ( .A(Reg_data[347]), .Y(register__net106155) );
  BUFx4f_ASAP7_75t_R register___U11327 ( .A(register__net97117), .Y(register__net106156) );
  BUFx4f_ASAP7_75t_R register___U11328 ( .A(register__net97117), .Y(register__net106157) );
  BUFx4f_ASAP7_75t_R register___U11329 ( .A(register__net106154), .Y(register__net97118) );
  BUFx3_ASAP7_75t_R register___U11330 ( .A(register__net106030), .Y(register__net106029) );
  BUFx2_ASAP7_75t_R register___U11331 ( .A(Reg_data[953]), .Y(register__net106030) );
  BUFx12f_ASAP7_75t_R register___U11332 ( .A(register__net88473), .Y(register__net88472) );
  BUFx3_ASAP7_75t_R register___U11333 ( .A(register__n7398), .Y(register__n7397) );
  BUFx2_ASAP7_75t_R register___U11334 ( .A(Reg_data[949]), .Y(register__n7398) );
  BUFx3_ASAP7_75t_R register___U11335 ( .A(register__n9581), .Y(register__n7399) );
  BUFx2_ASAP7_75t_R register___U11336 ( .A(register__n9581), .Y(register__n7400) );
  BUFx4f_ASAP7_75t_R register___U11337 ( .A(register__n9581), .Y(register__n7401) );
  BUFx3_ASAP7_75t_R register___U11338 ( .A(register__n7403), .Y(register__n7402) );
  BUFx2_ASAP7_75t_R register___U11339 ( .A(Reg_data[930]), .Y(register__n7403) );
  BUFx3_ASAP7_75t_R register___U11340 ( .A(register__n7405), .Y(register__n7404) );
  BUFx2_ASAP7_75t_R register___U11341 ( .A(Reg_data[916]), .Y(register__n7405) );
  BUFx3_ASAP7_75t_R register___U11342 ( .A(register__n7407), .Y(register__n7406) );
  BUFx2_ASAP7_75t_R register___U11343 ( .A(Reg_data[912]), .Y(register__n7407) );
  BUFx3_ASAP7_75t_R register___U11344 ( .A(register__n7409), .Y(register__n7408) );
  BUFx2_ASAP7_75t_R register___U11345 ( .A(Reg_data[897]), .Y(register__n7409) );
  BUFx3_ASAP7_75t_R register___U11346 ( .A(register__n7411), .Y(register__n7410) );
  BUFx2_ASAP7_75t_R register___U11347 ( .A(Reg_data[724]), .Y(register__n7411) );
  BUFx3_ASAP7_75t_R register___U11348 ( .A(register__n7413), .Y(register__n7412) );
  BUFx2_ASAP7_75t_R register___U11349 ( .A(Reg_data[722]), .Y(register__n7413) );
  BUFx3_ASAP7_75t_R register___U11350 ( .A(register__net105992), .Y(register__net105991) );
  BUFx2_ASAP7_75t_R register___U11351 ( .A(Reg_data[633]), .Y(register__net105992) );
  BUFx3_ASAP7_75t_R register___U11352 ( .A(register__n7415), .Y(register__n7414) );
  BUFx2_ASAP7_75t_R register___U11353 ( .A(Reg_data[630]), .Y(register__n7415) );
  BUFx3_ASAP7_75t_R register___U11354 ( .A(register__n7417), .Y(register__n7416) );
  BUFx2_ASAP7_75t_R register___U11355 ( .A(Reg_data[629]), .Y(register__n7417) );
  BUFx3_ASAP7_75t_R register___U11356 ( .A(register__n7419), .Y(register__n7418) );
  BUFx2_ASAP7_75t_R register___U11357 ( .A(Reg_data[624]), .Y(register__n7419) );
  BUFx3_ASAP7_75t_R register___U11358 ( .A(register__n7421), .Y(register__n7420) );
  BUFx2_ASAP7_75t_R register___U11359 ( .A(Reg_data[566]), .Y(register__n7421) );
  BUFx3_ASAP7_75t_R register___U11360 ( .A(register__n7423), .Y(register__n7422) );
  BUFx2_ASAP7_75t_R register___U11361 ( .A(Reg_data[552]), .Y(register__n7423) );
  BUFx3_ASAP7_75t_R register___U11362 ( .A(register__n7425), .Y(register__n7424) );
  BUFx2_ASAP7_75t_R register___U11363 ( .A(Reg_data[548]), .Y(register__n7425) );
  BUFx3_ASAP7_75t_R register___U11364 ( .A(register__n7427), .Y(register__n7426) );
  BUFx2_ASAP7_75t_R register___U11365 ( .A(Reg_data[547]), .Y(register__n7427) );
  BUFx3_ASAP7_75t_R register___U11366 ( .A(register__n7429), .Y(register__n7428) );
  BUFx2_ASAP7_75t_R register___U11367 ( .A(Reg_data[545]), .Y(register__n7429) );
  BUFx3_ASAP7_75t_R register___U11368 ( .A(register__n7431), .Y(register__n7430) );
  BUFx2_ASAP7_75t_R register___U11369 ( .A(Reg_data[512]), .Y(register__n7431) );
  BUFx3_ASAP7_75t_R register___U11370 ( .A(register__n7433), .Y(register__n7432) );
  BUFx2_ASAP7_75t_R register___U11371 ( .A(Reg_data[468]), .Y(register__n7433) );
  BUFx3_ASAP7_75t_R register___U11372 ( .A(register__n7435), .Y(register__n7434) );
  BUFx2_ASAP7_75t_R register___U11373 ( .A(Reg_data[466]), .Y(register__n7435) );
  BUFx3_ASAP7_75t_R register___U11374 ( .A(register__n10489), .Y(register__n7436) );
  BUFx2_ASAP7_75t_R register___U11375 ( .A(register__n10489), .Y(register__n7437) );
  BUFx4f_ASAP7_75t_R register___U11376 ( .A(register__n10489), .Y(register__n7438) );
  BUFx3_ASAP7_75t_R register___U11377 ( .A(register__n7440), .Y(register__n7439) );
  BUFx2_ASAP7_75t_R register___U11378 ( .A(Reg_data[464]), .Y(register__n7440) );
  BUFx3_ASAP7_75t_R register___U11379 ( .A(register__n7442), .Y(register__n7441) );
  BUFx2_ASAP7_75t_R register___U11380 ( .A(Reg_data[352]), .Y(register__n7442) );
  BUFx3_ASAP7_75t_R register___U11381 ( .A(register__n7444), .Y(register__n7443) );
  BUFx2_ASAP7_75t_R register___U11382 ( .A(Reg_data[342]), .Y(register__n7444) );
  BUFx3_ASAP7_75t_R register___U11383 ( .A(register__n7446), .Y(register__n7445) );
  BUFx2_ASAP7_75t_R register___U11384 ( .A(Reg_data[296]), .Y(register__n7446) );
  BUFx3_ASAP7_75t_R register___U11385 ( .A(register__net105922), .Y(register__net105921) );
  BUFx2_ASAP7_75t_R register___U11386 ( .A(Reg_data[294]), .Y(register__net105922) );
  BUFx3_ASAP7_75t_R register___U11387 ( .A(register__n7448), .Y(register__n7447) );
  BUFx2_ASAP7_75t_R register___U11388 ( .A(Reg_data[182]), .Y(register__n7448) );
  BUFx3_ASAP7_75t_R register___U11389 ( .A(register__net105914), .Y(register__net105913) );
  BUFx2_ASAP7_75t_R register___U11390 ( .A(Reg_data[165]), .Y(register__net105914) );
  BUFx3_ASAP7_75t_R register___U11391 ( .A(register__net105910), .Y(register__net105909) );
  BUFx2_ASAP7_75t_R register___U11392 ( .A(Reg_data[89]), .Y(register__net105910) );
  BUFx3_ASAP7_75t_R register___U11393 ( .A(register__n7450), .Y(register__n7449) );
  BUFx2_ASAP7_75t_R register___U11394 ( .A(Reg_data[68]), .Y(register__n7450) );
  BUFx3_ASAP7_75t_R register___U11395 ( .A(register__n7452), .Y(register__n7451) );
  BUFx2_ASAP7_75t_R register___U11396 ( .A(Reg_data[867]), .Y(register__n7452) );
  BUFx3_ASAP7_75t_R register___U11397 ( .A(register__n7454), .Y(register__n7453) );
  BUFx2_ASAP7_75t_R register___U11398 ( .A(Reg_data[214]), .Y(register__n7454) );
  BUFx3_ASAP7_75t_R register___U11399 ( .A(register__n7456), .Y(register__n7455) );
  BUFx2_ASAP7_75t_R register___U11400 ( .A(Reg_data[213]), .Y(register__n7456) );
  BUFx2_ASAP7_75t_R register___U11401 ( .A(register__n10054), .Y(register__n7457) );
  BUFx2_ASAP7_75t_R register___U11402 ( .A(register__n10054), .Y(register__n7458) );
  BUFx4f_ASAP7_75t_R register___U11403 ( .A(register__n10054), .Y(register__n7459) );
  BUFx3_ASAP7_75t_R register___U11404 ( .A(register__net105884), .Y(register__net105883) );
  BUFx2_ASAP7_75t_R register___U11405 ( .A(Reg_data[198]), .Y(register__net105884) );
  BUFx3_ASAP7_75t_R register___U11406 ( .A(register__net105880), .Y(register__net105879) );
  BUFx2_ASAP7_75t_R register___U11407 ( .A(Reg_data[197]), .Y(register__net105880) );
  BUFx3_ASAP7_75t_R register___U11408 ( .A(register__n7461), .Y(register__n7460) );
  BUFx2_ASAP7_75t_R register___U11409 ( .A(Reg_data[196]), .Y(register__n7461) );
  BUFx3_ASAP7_75t_R register___U11410 ( .A(register__n7463), .Y(register__n7462) );
  BUFx2_ASAP7_75t_R register___U11411 ( .A(Reg_data[195]), .Y(register__n7463) );
  BUFx3_ASAP7_75t_R register___U11412 ( .A(register__n7465), .Y(register__n7464) );
  BUFx2_ASAP7_75t_R register___U11413 ( .A(Reg_data[193]), .Y(register__n7465) );
  BUFx4f_ASAP7_75t_R register___U11414 ( .A(register__n8791), .Y(register__n7466) );
  BUFx2_ASAP7_75t_R register___U11415 ( .A(register__n8791), .Y(register__n7467) );
  BUFx3_ASAP7_75t_R register___U11416 ( .A(register__n8791), .Y(register__n7468) );
  BUFx3_ASAP7_75t_R register___U11417 ( .A(register__n7470), .Y(register__n7469) );
  BUFx2_ASAP7_75t_R register___U11418 ( .A(Reg_data[20]), .Y(register__n7470) );
  BUFx3_ASAP7_75t_R register___U11419 ( .A(register__n7472), .Y(register__n7471) );
  BUFx2_ASAP7_75t_R register___U11420 ( .A(Reg_data[18]), .Y(register__n7472) );
  BUFx3_ASAP7_75t_R register___U11421 ( .A(register__n7474), .Y(register__n7473) );
  BUFx2_ASAP7_75t_R register___U11422 ( .A(Reg_data[200]), .Y(register__n7474) );
  BUFx3_ASAP7_75t_R register___U11423 ( .A(register__n7476), .Y(register__n7475) );
  BUFx2_ASAP7_75t_R register___U11424 ( .A(Reg_data[224]), .Y(register__n7476) );
  BUFx2_ASAP7_75t_R register___U11425 ( .A(register__n10070), .Y(register__n7477) );
  BUFx2_ASAP7_75t_R register___U11426 ( .A(register__n10070), .Y(register__n7478) );
  BUFx4f_ASAP7_75t_R register___U11427 ( .A(register__n10070), .Y(register__n7479) );
  BUFx3_ASAP7_75t_R register___U11428 ( .A(register__n7481), .Y(register__n7480) );
  BUFx2_ASAP7_75t_R register___U11429 ( .A(Reg_data[33]), .Y(register__n7481) );
  BUFx3_ASAP7_75t_R register___U11430 ( .A(register__n7483), .Y(register__n7482) );
  BUFx2_ASAP7_75t_R register___U11431 ( .A(Reg_data[35]), .Y(register__n7483) );
  BUFx3_ASAP7_75t_R register___U11432 ( .A(register__n7485), .Y(register__n7484) );
  BUFx2_ASAP7_75t_R register___U11433 ( .A(Reg_data[244]), .Y(register__n7485) );
  BUFx2_ASAP7_75t_R register___U11434 ( .A(register__n10086), .Y(register__n7487) );
  BUFx4f_ASAP7_75t_R register___U11435 ( .A(register__n10086), .Y(register__n7488) );
  BUFx3_ASAP7_75t_R register___U11436 ( .A(register__n7490), .Y(register__n7489) );
  BUFx2_ASAP7_75t_R register___U11437 ( .A(Reg_data[240]), .Y(register__n7490) );
  BUFx4f_ASAP7_75t_R register___U11438 ( .A(register__net123812), .Y(register__net105809) );
  BUFx2_ASAP7_75t_R register___U11439 ( .A(Reg_data[939]), .Y(register__net105810) );
  BUFx12f_ASAP7_75t_R register___U11440 ( .A(register__net90718), .Y(register__net90717) );
  BUFx6f_ASAP7_75t_R register___U11441 ( .A(register__net105809), .Y(register__net90718) );
  BUFx3_ASAP7_75t_R register___U11442 ( .A(register__n7492), .Y(register__n7491) );
  BUFx2_ASAP7_75t_R register___U11443 ( .A(Reg_data[301]), .Y(register__n7492) );
  BUFx3_ASAP7_75t_R register___U11444 ( .A(register__net105802), .Y(register__net105801) );
  BUFx2_ASAP7_75t_R register___U11445 ( .A(Reg_data[11]), .Y(register__net105802) );
  BUFx3_ASAP7_75t_R register___U11446 ( .A(register__net105795), .Y(register__net105794) );
  BUFx2_ASAP7_75t_R register___U11447 ( .A(Reg_data[299]), .Y(register__net105795) );
  BUFx12f_ASAP7_75t_R register___U11448 ( .A(register__net90674), .Y(register__net90673) );
  BUFx3_ASAP7_75t_R register___U11449 ( .A(register__net105791), .Y(register__net105790) );
  BUFx2_ASAP7_75t_R register___U11450 ( .A(Reg_data[427]), .Y(register__net105791) );
  BUFx3_ASAP7_75t_R register___U11451 ( .A(register__net105787), .Y(register__net105786) );
  BUFx2_ASAP7_75t_R register___U11452 ( .A(Reg_data[203]), .Y(register__net105787) );
  BUFx3_ASAP7_75t_R register___U11453 ( .A(register__net105783), .Y(register__net105782) );
  BUFx2_ASAP7_75t_R register___U11454 ( .A(Reg_data[655]), .Y(register__net105783) );
  BUFx3_ASAP7_75t_R register___U11455 ( .A(register__n7494), .Y(register__n7493) );
  BUFx2_ASAP7_75t_R register___U11456 ( .A(Reg_data[461]), .Y(register__n7494) );
  BUFx3_ASAP7_75t_R register___U11457 ( .A(register__n7496), .Y(register__n7495) );
  BUFx2_ASAP7_75t_R register___U11458 ( .A(Reg_data[909]), .Y(register__n7496) );
  BUFx3_ASAP7_75t_R register___U11459 ( .A(register__n7498), .Y(register__n7497) );
  BUFx2_ASAP7_75t_R register___U11460 ( .A(Reg_data[460]), .Y(register__n7498) );
  BUFx3_ASAP7_75t_R register___U11461 ( .A(register__n7500), .Y(register__n7499) );
  BUFx2_ASAP7_75t_R register___U11462 ( .A(Reg_data[366]), .Y(register__n7500) );
  BUFx3_ASAP7_75t_R register___U11463 ( .A(register__n7502), .Y(register__n7501) );
  BUFx2_ASAP7_75t_R register___U11464 ( .A(Reg_data[314]), .Y(register__n7502) );
  BUFx3_ASAP7_75t_R register___U11465 ( .A(register__n7504), .Y(register__n7503) );
  BUFx2_ASAP7_75t_R register___U11466 ( .A(Reg_data[300]), .Y(register__n7504) );
  BUFx3_ASAP7_75t_R register___U11467 ( .A(register__net105755), .Y(register__net105754) );
  BUFx2_ASAP7_75t_R register___U11468 ( .A(Reg_data[303]), .Y(register__net105755) );
  BUFx3_ASAP7_75t_R register___U11469 ( .A(register__n7506), .Y(register__n7505) );
  BUFx2_ASAP7_75t_R register___U11470 ( .A(Reg_data[841]), .Y(register__n7506) );
  BUFx3_ASAP7_75t_R register___U11471 ( .A(register__n7508), .Y(register__n7507) );
  BUFx2_ASAP7_75t_R register___U11472 ( .A(Reg_data[81]), .Y(register__n7508) );
  BUFx3_ASAP7_75t_R register___U11473 ( .A(register__n7510), .Y(register__n7509) );
  BUFx2_ASAP7_75t_R register___U11474 ( .A(Reg_data[220]), .Y(register__n7510) );
  BUFx3_ASAP7_75t_R register___U11475 ( .A(register__net105739), .Y(register__net105738) );
  BUFx2_ASAP7_75t_R register___U11476 ( .A(Reg_data[408]), .Y(register__net105739) );
  BUFx3_ASAP7_75t_R register___U11477 ( .A(register__net105735), .Y(register__net105734) );
  BUFx2_ASAP7_75t_R register___U11478 ( .A(Reg_data[56]), .Y(register__net105735) );
  BUFx3_ASAP7_75t_R register___U11479 ( .A(register__n7512), .Y(register__n7511) );
  BUFx2_ASAP7_75t_R register___U11480 ( .A(Reg_data[903]), .Y(register__n7512) );
  BUFx4f_ASAP7_75t_R register___U11481 ( .A(register__n9782), .Y(register__n7513) );
  BUFx2_ASAP7_75t_R register___U11482 ( .A(register__n9782), .Y(register__n7514) );
  BUFx3_ASAP7_75t_R register___U11483 ( .A(register__n9782), .Y(register__n7515) );
  BUFx3_ASAP7_75t_R register___U11484 ( .A(register__n7517), .Y(register__n7516) );
  BUFx2_ASAP7_75t_R register___U11485 ( .A(Reg_data[158]), .Y(register__n7517) );
  BUFx3_ASAP7_75t_R register___U11486 ( .A(register__n7519), .Y(register__n7518) );
  BUFx2_ASAP7_75t_R register___U11487 ( .A(Reg_data[412]), .Y(register__n7519) );
  BUFx2_ASAP7_75t_R register___U11488 ( .A(register__n9808), .Y(register__n7520) );
  BUFx2_ASAP7_75t_R register___U11489 ( .A(register__n9808), .Y(register__n7521) );
  BUFx4f_ASAP7_75t_R register___U11490 ( .A(register__n9808), .Y(register__n7522) );
  BUFx3_ASAP7_75t_R register___U11491 ( .A(register__n7524), .Y(register__n7523) );
  BUFx2_ASAP7_75t_R register___U11492 ( .A(Reg_data[508]), .Y(register__n7524) );
  BUFx3_ASAP7_75t_R register___U11493 ( .A(register__n7526), .Y(register__n7525) );
  BUFx2_ASAP7_75t_R register___U11494 ( .A(Reg_data[908]), .Y(register__n7526) );
  BUFx3_ASAP7_75t_R register___U11495 ( .A(register__n7528), .Y(register__n7527) );
  BUFx2_ASAP7_75t_R register___U11496 ( .A(Reg_data[684]), .Y(register__n7528) );
  BUFx3_ASAP7_75t_R register___U11497 ( .A(register__n7530), .Y(register__n7529) );
  BUFx2_ASAP7_75t_R register___U11498 ( .A(Reg_data[83]), .Y(register__n7530) );
  BUFx3_ASAP7_75t_R register___U11499 ( .A(register__n7532), .Y(register__n7531) );
  BUFx2_ASAP7_75t_R register___U11500 ( .A(Reg_data[691]), .Y(register__n7532) );
  BUFx3_ASAP7_75t_R register___U11501 ( .A(register__net105687), .Y(register__net105686) );
  BUFx2_ASAP7_75t_R register___U11502 ( .A(Reg_data[362]), .Y(register__net105687) );
  BUFx3_ASAP7_75t_R register___U11503 ( .A(register__net105683), .Y(register__net105682) );
  BUFx2_ASAP7_75t_R register___U11504 ( .A(Reg_data[458]), .Y(register__net105683) );
  BUFx3_ASAP7_75t_R register___U11505 ( .A(register__net105679), .Y(register__net105678) );
  BUFx2_ASAP7_75t_R register___U11506 ( .A(Reg_data[10]), .Y(register__net105679) );
  BUFx4f_ASAP7_75t_R register___U11507 ( .A(register__n5177), .Y(register__n7533) );
  BUFx2_ASAP7_75t_R register___U11508 ( .A(Reg_data[951]), .Y(register__n7534) );
  BUFx12f_ASAP7_75t_R register___U11509 ( .A(register__n9837), .Y(register__n7535) );
  BUFx12f_ASAP7_75t_R register___U11510 ( .A(register__n7535), .Y(register__n9836) );
  BUFx6f_ASAP7_75t_R register___U11511 ( .A(register__n7533), .Y(register__n9837) );
  BUFx3_ASAP7_75t_R register___U11512 ( .A(register__n7537), .Y(register__n7536) );
  BUFx2_ASAP7_75t_R register___U11513 ( .A(Reg_data[891]), .Y(register__n7537) );
  BUFx4f_ASAP7_75t_R register___U11514 ( .A(register__n9838), .Y(register__n7538) );
  BUFx2_ASAP7_75t_R register___U11515 ( .A(register__n9838), .Y(register__n7539) );
  BUFx2_ASAP7_75t_R register___U11516 ( .A(register__n9838), .Y(register__n7540) );
  BUFx3_ASAP7_75t_R register___U11517 ( .A(register__n7542), .Y(register__n7541) );
  BUFx2_ASAP7_75t_R register___U11518 ( .A(Reg_data[201]), .Y(register__n7542) );
  BUFx3_ASAP7_75t_R register___U11519 ( .A(register__n7544), .Y(register__n7543) );
  BUFx2_ASAP7_75t_R register___U11520 ( .A(Reg_data[9]), .Y(register__n7544) );
  BUFx3_ASAP7_75t_R register___U11521 ( .A(register__n7546), .Y(register__n7545) );
  BUFx2_ASAP7_75t_R register___U11522 ( .A(Reg_data[538]), .Y(register__n7546) );
  BUFx3_ASAP7_75t_R register___U11523 ( .A(register__n7548), .Y(register__n7547) );
  BUFx2_ASAP7_75t_R register___U11524 ( .A(Reg_data[927]), .Y(register__n7548) );
  BUFx2_ASAP7_75t_R register___U11525 ( .A(register__n9859), .Y(register__n7549) );
  BUFx2_ASAP7_75t_R register___U11526 ( .A(register__n9859), .Y(register__n7550) );
  BUFx4f_ASAP7_75t_R register___U11527 ( .A(register__n9859), .Y(register__n7551) );
  BUFx3_ASAP7_75t_R register___U11528 ( .A(register__n7553), .Y(register__n7552) );
  BUFx2_ASAP7_75t_R register___U11529 ( .A(Reg_data[937]), .Y(register__n7553) );
  BUFx3_ASAP7_75t_R register___U11530 ( .A(register__n9865), .Y(register__n7554) );
  BUFx2_ASAP7_75t_R register___U11531 ( .A(register__n9865), .Y(register__n7555) );
  BUFx4f_ASAP7_75t_R register___U11532 ( .A(register__n9865), .Y(register__n7556) );
  BUFx3_ASAP7_75t_R register___U11533 ( .A(register__n7558), .Y(register__n7557) );
  BUFx2_ASAP7_75t_R register___U11534 ( .A(Reg_data[90]), .Y(register__n7558) );
  BUFx3_ASAP7_75t_R register___U11535 ( .A(register__n7560), .Y(register__n7559) );
  BUFx2_ASAP7_75t_R register___U11536 ( .A(Reg_data[529]), .Y(register__n7560) );
  BUFx2_ASAP7_75t_R register___U11537 ( .A(register__n10309), .Y(register__n7561) );
  BUFx2_ASAP7_75t_R register___U11538 ( .A(register__n10309), .Y(register__n7562) );
  BUFx4f_ASAP7_75t_R register___U11539 ( .A(register__n10309), .Y(register__n7563) );
  BUFx4f_ASAP7_75t_R register___U11540 ( .A(register__n7134), .Y(register__n7564) );
  BUFx2_ASAP7_75t_R register___U11541 ( .A(Reg_data[721]), .Y(register__n7565) );
  BUFx12f_ASAP7_75t_R register___U11542 ( .A(register__n10318), .Y(register__n7566) );
  BUFx12f_ASAP7_75t_R register___U11543 ( .A(register__n7566), .Y(register__n10317) );
  BUFx6f_ASAP7_75t_R register___U11544 ( .A(register__n7564), .Y(register__n10318) );
  BUFx3_ASAP7_75t_R register___U11545 ( .A(register__n7568), .Y(register__n7567) );
  BUFx2_ASAP7_75t_R register___U11546 ( .A(Reg_data[475]), .Y(register__n7568) );
  BUFx2_ASAP7_75t_R register___U11547 ( .A(Reg_data[59]), .Y(register__n7570) );
  BUFx3_ASAP7_75t_R register___U11548 ( .A(register__n7572), .Y(register__n7571) );
  BUFx2_ASAP7_75t_R register___U11549 ( .A(Reg_data[383]), .Y(register__n7572) );
  BUFx2_ASAP7_75t_R register___U11550 ( .A(register__n9893), .Y(register__n7573) );
  BUFx6f_ASAP7_75t_R register___U11551 ( .A(register__n9893), .Y(register__n7574) );
  BUFx3_ASAP7_75t_R register___U11552 ( .A(register__net105583), .Y(register__net105582) );
  BUFx2_ASAP7_75t_R register___U11553 ( .A(Reg_data[477]), .Y(register__net105583) );
  BUFx2_ASAP7_75t_R register___U11554 ( .A(Reg_data[637]), .Y(register__net105576) );
  BUFx4f_ASAP7_75t_R register___U11555 ( .A(register__n11459), .Y(register__n7575) );
  INVx2_ASAP7_75t_R register___U11556 ( .A(register__n7148), .Y(register__n11459) );
  BUFx6f_ASAP7_75t_R register___U11557 ( .A(register__n8333), .Y(register__n8332) );
  BUFx4f_ASAP7_75t_R register___U11558 ( .A(register__n9217), .Y(register__n11708) );
  INVx1_ASAP7_75t_R register___U11559 ( .A(register__n11708), .Y(register__n7576) );
  BUFx6f_ASAP7_75t_R register___U11560 ( .A(register__n9218), .Y(register__n9217) );
  BUFx4f_ASAP7_75t_R register___U11561 ( .A(register__n11022), .Y(register__n7577) );
  INVx2_ASAP7_75t_R register___U11562 ( .A(register__n6824), .Y(register__n11022) );
  BUFx6f_ASAP7_75t_R register___U11563 ( .A(register__n8739), .Y(register__n8738) );
  BUFx4f_ASAP7_75t_R register___U11564 ( .A(register__n11374), .Y(register__n7578) );
  INVx2_ASAP7_75t_R register___U11565 ( .A(register__n8740), .Y(register__n11374) );
  BUFx6f_ASAP7_75t_R register___U11566 ( .A(register__n8741), .Y(register__n8740) );
  BUFx4f_ASAP7_75t_R register___U11567 ( .A(register__n11481), .Y(register__n7579) );
  INVx2_ASAP7_75t_R register___U11568 ( .A(register__n7984), .Y(register__n11481) );
  BUFx6f_ASAP7_75t_R register___U11569 ( .A(register__n7985), .Y(register__n7984) );
  INVx2_ASAP7_75t_R register___U11570 ( .A(register__n8706), .Y(register__n10533) );
  BUFx6f_ASAP7_75t_R register___U11571 ( .A(register__n8707), .Y(register__n8706) );
  BUFx4f_ASAP7_75t_R register___U11572 ( .A(register__n10937), .Y(register__n7581) );
  INVx2_ASAP7_75t_R register___U11573 ( .A(register__n7982), .Y(register__n10937) );
  BUFx6f_ASAP7_75t_R register___U11574 ( .A(register__n7983), .Y(register__n7982) );
  INVx2_ASAP7_75t_R register___U11575 ( .A(register__net102363), .Y(register__net105530) );
  BUFx6f_ASAP7_75t_R register___U11576 ( .A(register__net102364), .Y(register__net102363) );
  BUFx6f_ASAP7_75t_R register___U11577 ( .A(register__net97186), .Y(register__net97185) );
  BUFx4f_ASAP7_75t_R register___U11578 ( .A(register__n10683), .Y(register__n7582) );
  INVx2_ASAP7_75t_R register___U11579 ( .A(register__n8736), .Y(register__n10683) );
  BUFx6f_ASAP7_75t_R register___U11580 ( .A(register__n8737), .Y(register__n8736) );
  BUFx6f_ASAP7_75t_R register___U11581 ( .A(register__net102360), .Y(register__net102359) );
  BUFx4f_ASAP7_75t_R register___U11582 ( .A(register__n10891), .Y(register__n7583) );
  INVx2_ASAP7_75t_R register___U11583 ( .A(register__n8732), .Y(register__n10891) );
  BUFx6f_ASAP7_75t_R register___U11584 ( .A(register__n8733), .Y(register__n8732) );
  BUFx3_ASAP7_75t_R register___U11585 ( .A(register__n11413), .Y(register__n7584) );
  BUFx2_ASAP7_75t_R register___U11586 ( .A(register__n11413), .Y(register__n7585) );
  INVx2_ASAP7_75t_R register___U11587 ( .A(register__n8728), .Y(register__n11413) );
  BUFx6f_ASAP7_75t_R register___U11588 ( .A(register__n8729), .Y(register__n8728) );
  INVx2_ASAP7_75t_R register___U11589 ( .A(register__net97237), .Y(register__net105496) );
  BUFx6f_ASAP7_75t_R register___U11590 ( .A(register__net97238), .Y(register__net97237) );
  BUFx4f_ASAP7_75t_R register___U11591 ( .A(register__n11246), .Y(register__n7586) );
  INVx2_ASAP7_75t_R register___U11592 ( .A(register__n8712), .Y(register__n11246) );
  BUFx6f_ASAP7_75t_R register___U11593 ( .A(register__n8713), .Y(register__n8712) );
  INVx2_ASAP7_75t_R register___U11594 ( .A(register__net94144), .Y(register__net105488) );
  BUFx6f_ASAP7_75t_R register___U11595 ( .A(register__net94145), .Y(register__net94144) );
  OA22x2_ASAP7_75t_R register___U11596 ( .A1(register__n11996), .A2(register__n4267), .B1(register__n8912), .B2(register__n3479), 
        .Y(register__n12634) );
  INVx1_ASAP7_75t_R register___U11597 ( .A(register__n4509), .Y(register__n7587) );
  OA22x2_ASAP7_75t_R register___U11598 ( .A1(register__n12261), .A2(register__n4267), .B1(register__n8931), .B2(register__n11902), 
        .Y(register__n12618) );
  INVx1_ASAP7_75t_R register___U11599 ( .A(register__n4005), .Y(register__n7588) );
  OA22x2_ASAP7_75t_R register___U11600 ( .A1(register__net64942), .A2(register__n4267), .B1(register__n9714), .B2(
        n11824), .Y(register__n12632) );
  INVx1_ASAP7_75t_R register___U11601 ( .A(register__n4513), .Y(register__n7589) );
  OA22x2_ASAP7_75t_R register___U11602 ( .A1(register__net63180), .A2(register__n1989), .B1(register__net89741), .B2(
        n4952), .Y(register__n13339) );
  INVx1_ASAP7_75t_R register___U11603 ( .A(register__n3897), .Y(register__n7590) );
  OA22x2_ASAP7_75t_R register___U11604 ( .A1(register__n12254), .A2(register__n1988), .B1(register__n10080), .B2(register__n4373), 
        .Y(register__n13345) );
  OA22x2_ASAP7_75t_R register___U11605 ( .A1(register__n12092), .A2(register__n4267), .B1(register__n9774), .B2(register__n11821), 
        .Y(register__n12627) );
  OA22x2_ASAP7_75t_R register___U11606 ( .A1(register__net64690), .A2(register__n4267), .B1(register__n9780), .B2(register__n3756), .Y(register__n12629) );
  INVx1_ASAP7_75t_R register___U11607 ( .A(register__n4415), .Y(register__n7591) );
  OA22x2_ASAP7_75t_R register___U11608 ( .A1(register__net63264), .A2(register__n11900), .B1(register__net90257), .B2(
        n3263), .Y(register__n12612) );
  OA22x2_ASAP7_75t_R register___U11609 ( .A1(register__n12192), .A2(register__n1989), .B1(register__n10462), .B2(register__n6721), 
        .Y(register__n13347) );
  INVx2_ASAP7_75t_R register___U11610 ( .A(register__net91940), .Y(register__net64442) );
  OA22x2_ASAP7_75t_R register___U11611 ( .A1(register__net62674), .A2(register__n11900), .B1(register__n9857), .B2(
        n1510), .Y(register__n12606) );
  INVx1_ASAP7_75t_R register___U11612 ( .A(register__n4367), .Y(register__n7594) );
  INVx1_ASAP7_75t_R register___U11613 ( .A(register__n4369), .Y(register__n7595) );
  INVx1_ASAP7_75t_R register___U11614 ( .A(register__n5110), .Y(register__n7597) );
  INVx1_ASAP7_75t_R register___U11615 ( .A(register__n5560), .Y(register__n7600) );
  INVx1_ASAP7_75t_R register___U11616 ( .A(register__n10690), .Y(register__n7602) );
  INVx1_ASAP7_75t_R register___U11617 ( .A(register__n5299), .Y(register__n7608) );
  BUFx12f_ASAP7_75t_R register___U11618 ( .A(register__n11980), .Y(register__n7609) );
  BUFx6f_ASAP7_75t_R register___U11619 ( .A(register__n11972), .Y(register__n11976) );
  BUFx6f_ASAP7_75t_R register___U11620 ( .A(register__n3833), .Y(register__n11977) );
  OA22x2_ASAP7_75t_R register___U11621 ( .A1(register__n12376), .A2(register__n4267), .B1(register__n7703), .B2(register__n3547), 
        .Y(register__n12614) );
  OA22x2_ASAP7_75t_R register___U11622 ( .A1(register__net64668), .A2(register__n1735), .B1(register__n8132), .B2(register__n3352), .Y(register__n13257) );
  BUFx6f_ASAP7_75t_R register___U11623 ( .A(register__net64816), .Y(register__net64800) );
  BUFx6f_ASAP7_75t_R register___U11624 ( .A(register__net64796), .Y(register__net64808) );
  OA22x2_ASAP7_75t_R register___U11625 ( .A1(register__n12321), .A2(register__n188), .B1(register__n9611), .B2(register__n215), 
        .Y(register__n12672) );
  INVx1_ASAP7_75t_R register___U11626 ( .A(register__n7116), .Y(register__n7615) );
  OA22x2_ASAP7_75t_R register___U11627 ( .A1(register__n12051), .A2(register__n1988), .B1(register__n10463), .B2(register__n11850), .Y(register__n13353) );
  OA22x2_ASAP7_75t_R register___U11628 ( .A1(register__net64344), .A2(register__n4033), .B1(register__net93817), .B2(
        n3384), .Y(register__n12541) );
  OA22x2_ASAP7_75t_R register___U11629 ( .A1(register__net62672), .A2(register__n196), .B1(register__n8781), .B2(register__n216), 
        .Y(register__n12661) );
  OA22x2_ASAP7_75t_R register___U11630 ( .A1(register__net64844), .A2(register__n3991), .B1(register__net93837), .B2(
        n4034), .Y(register__n12547) );
  INVx1_ASAP7_75t_R register___U11631 ( .A(register__n12547), .Y(register__n7619) );
  OA22x2_ASAP7_75t_R register___U11632 ( .A1(register__n11995), .A2(register__n190), .B1(register__n9617), .B2(register__n209), 
        .Y(register__n12689) );
  OA22x2_ASAP7_75t_R register___U11633 ( .A1(register__n12194), .A2(register__n1702), .B1(register__n10006), .B2(register__n1717), 
        .Y(register__n13249) );
  INVx1_ASAP7_75t_R register___U11634 ( .A(register__n4210), .Y(register__n7621) );
  OA22x2_ASAP7_75t_R register___U11635 ( .A1(register__net64920), .A2(register__n1736), .B1(register__n10010), .B2(
        n4575), .Y(register__n13260) );
  OA22x2_ASAP7_75t_R register___U11636 ( .A1(register__n11921), .A2(register__n1989), .B1(register__n10066), .B2(register__n2967), 
        .Y(register__n13357) );
  OA22x2_ASAP7_75t_R register___U11637 ( .A1(register__net129768), .A2(register__n4033), .B1(register__n9722), .B2(
        n4603), .Y(register__n12545) );
  INVx1_ASAP7_75t_R register___U11638 ( .A(register__n6504), .Y(register__n7622) );
  OA22x2_ASAP7_75t_R register___U11639 ( .A1(register__net63992), .A2(register__n4033), .B1(register__net93639), .B2(
        n11840), .Y(register__n12538) );
  INVx1_ASAP7_75t_R register___U11640 ( .A(register__n4430), .Y(register__n7623) );
  OA22x2_ASAP7_75t_R register___U11641 ( .A1(register__net64436), .A2(register__n184), .B1(register__net90649), .B2(
        n208), .Y(register__n12682) );
  INVx1_ASAP7_75t_R register___U11642 ( .A(register__n6787), .Y(register__n7624) );
  OA22x2_ASAP7_75t_R register___U11643 ( .A1(register__n12110), .A2(register__n1988), .B1(register__n10142), .B2(register__n5182), 
        .Y(register__n13350) );
  OA22x2_ASAP7_75t_R register___U11644 ( .A1(register__n12122), .A2(register__n177), .B1(register__n9812), .B2(register__n208), 
        .Y(register__n12680) );
  INVx1_ASAP7_75t_R register___U11645 ( .A(register__n12680), .Y(register__n7627) );
  OA22x2_ASAP7_75t_R register___U11646 ( .A1(register__n11951), .A2(register__n1700), .B1(register__n4182), .B2(register__n1731), 
        .Y(register__n13262) );
  INVx1_ASAP7_75t_R register___U11647 ( .A(register__n4058), .Y(register__n7629) );
  INVx4_ASAP7_75t_R register___U11648 ( .A(register__n11972), .Y(register__n11951) );
  OA22x2_ASAP7_75t_R register___U11649 ( .A1(register__net63344), .A2(register__n179), .B1(register__n8769), .B2(register__n210), 
        .Y(register__n12669) );
  INVx1_ASAP7_75t_R register___U11650 ( .A(register__n6783), .Y(register__n7630) );
  OA22x2_ASAP7_75t_R register___U11651 ( .A1(register__net63160), .A2(register__n4033), .B1(register__net93853), .B2(
        n11919), .Y(register__n12528) );
  INVx1_ASAP7_75t_R register___U11652 ( .A(register__n5747), .Y(register__n7631) );
  OA22x2_ASAP7_75t_R register___U11653 ( .A1(register__net63176), .A2(register__n191), .B1(register__net91021), .B2(
        n212), .Y(register__n12667) );
  OA22x2_ASAP7_75t_R register___U11654 ( .A1(register__net62648), .A2(register__n1988), .B1(register__n10325), .B2(
        n11732), .Y(register__n13335) );
  INVx5_ASAP7_75t_R register___U11655 ( .A(register__net62682), .Y(register__net62648) );
  INVx1_ASAP7_75t_R register___U11656 ( .A(register__n3030), .Y(register__n7634) );
  INVx1_ASAP7_75t_R register___U11657 ( .A(register__n3084), .Y(register__n7635) );
  INVx1_ASAP7_75t_R register___U11658 ( .A(register__n3086), .Y(register__n7636) );
  INVx1_ASAP7_75t_R register___U11659 ( .A(register__n3089), .Y(register__n7637) );
  INVx1_ASAP7_75t_R register___U11660 ( .A(register__n10857), .Y(register__n7640) );
  AO22x1_ASAP7_75t_R register___U11661 ( .A1(register__n7992), .A2(register__C6423_net61318), .B1(register__n10307), 
        .B2(register__n1442), .Y(register__n11462) );
  INVx1_ASAP7_75t_R register___U11662 ( .A(register__n11462), .Y(register__n7641) );
  INVx1_ASAP7_75t_R register___U11663 ( .A(register__n4329), .Y(register__n7642) );
  INVx1_ASAP7_75t_R register___U11664 ( .A(register__n10625), .Y(register__n7644) );
  INVx1_ASAP7_75t_R register___U11665 ( .A(register__n4247), .Y(register__n7645) );
  INVx1_ASAP7_75t_R register___U11666 ( .A(register__n10899), .Y(register__n7646) );
  INVx1_ASAP7_75t_R register___U11667 ( .A(register__n4250), .Y(register__n7647) );
  INVx1_ASAP7_75t_R register___U11668 ( .A(register__n4565), .Y(register__n7648) );
  INVx1_ASAP7_75t_R register___U11669 ( .A(register__n4566), .Y(register__n7649) );
  INVx1_ASAP7_75t_R register___U11670 ( .A(register__n4568), .Y(register__n7650) );
  INVx1_ASAP7_75t_R register___U11671 ( .A(register__n3182), .Y(register__n7651) );
  INVx1_ASAP7_75t_R register___U11672 ( .A(register__n3112), .Y(register__n7653) );
  BUFx6f_ASAP7_75t_R register___U11673 ( .A(register__net63044), .Y(register__net63018) );
  OA22x2_ASAP7_75t_R register___U11674 ( .A1(register__n6679), .A2(register__n4033), .B1(register__n9272), .B2(register__n4604), 
        .Y(register__n12534) );
  INVx1_ASAP7_75t_R register___U11675 ( .A(register__n4216), .Y(register__n7654) );
  OA22x2_ASAP7_75t_R register___U11676 ( .A1(register__net62840), .A2(register__n191), .B1(register__net96843), .B2(
        n220), .Y(register__n12663) );
  INVx1_ASAP7_75t_R register___U11677 ( .A(register__n12663), .Y(register__n7655) );
  BUFx12f_ASAP7_75t_R register___U11678 ( .A(register__n3217), .Y(register__n11806) );
  INVx1_ASAP7_75t_R register___U11679 ( .A(register__n6775), .Y(register__n7657) );
  BUFx2_ASAP7_75t_R register___U11680 ( .A(Reg_data[790]), .Y(register__n7658) );
  BUFx3_ASAP7_75t_R register___U11681 ( .A(register__n7658), .Y(register__n10956) );
  BUFx2_ASAP7_75t_R register___U11682 ( .A(Reg_data[783]), .Y(register__net104916) );
  BUFx3_ASAP7_75t_R register___U11683 ( .A(register__net104916), .Y(register__C6423_net60878) );
  OR3x1_ASAP7_75t_R register___U11684 ( .A(register__n5328), .B(register__n7666), .C(register__n7664), .Y(register__n11322) );
  OA22x2_ASAP7_75t_R register___U11685 ( .A1(register__net131654), .A2(register__n8001), .B1(register__net130175), .B2(
        n8359), .Y(register__n11325) );
  INVx1_ASAP7_75t_R register___U11686 ( .A(register__n5324), .Y(register__n7664) );
  INVx1_ASAP7_75t_R register___U11687 ( .A(register__n5326), .Y(register__n7665) );
  OA22x2_ASAP7_75t_R register___U11688 ( .A1(register__n713), .A2(register__n7247), .B1(register__n353), .B2(register__n6984), 
        .Y(register__n11324) );
  INVx1_ASAP7_75t_R register___U11689 ( .A(register__n5329), .Y(register__n7666) );
  OR3x1_ASAP7_75t_R register___U11690 ( .A(register__n5038), .B(register__n7669), .C(register__n7667), .Y(register__n11263) );
  OA22x2_ASAP7_75t_R register___U11691 ( .A1(register__net131654), .A2(register__net101833), .B1(register__net130175), 
        .B2(register__net103300), .Y(register__n11265) );
  INVx1_ASAP7_75t_R register___U11692 ( .A(register__n5036), .Y(register__n7667) );
  OA22x2_ASAP7_75t_R register___U11693 ( .A1(register__n712), .A2(register__net107791), .B1(register__net149938), .B2(
        net109852), .Y(register__n11264) );
  INVx1_ASAP7_75t_R register___U11694 ( .A(register__n5039), .Y(register__n7669) );
  OR3x1_ASAP7_75t_R register___U11695 ( .A(register__n7), .B(register__n8), .C(register__register__n7671), .Y(register__n10550) );
  OA22x2_ASAP7_75t_R register___U11696 ( .A1(register__n420), .A2(register__n6488), .B1(register__n11180), .B2(register__n802), 
        .Y(register__n10553) );
  OA22x2_ASAP7_75t_R register___U11697 ( .A1(register__net107674), .A2(register__n5956), .B1(register__n1691), .B2(
        n7244), .Y(register__n10552) );
  OA22x2_ASAP7_75t_R register___U11698 ( .A1(register__net131654), .A2(register__n6483), .B1(register__net130175), .B2(
        n8587), .Y(register__n11433) );
  OA22x2_ASAP7_75t_R register___U11699 ( .A1(register__n710), .A2(register__n7093), .B1(register__n1114), .B2(register__n8216), 
        .Y(register__n11432) );
  INVx1_ASAP7_75t_R register___U11700 ( .A(register__n5121), .Y(register__n7673) );
  OA222x2_ASAP7_75t_R register___U11701 ( .A1(register__n1987), .A2(register__n10825), .B1(register__n1995), .B2(register__n10826), .C1(register__n1800), .C2(register__n6206), .Y(register__n11431) );
  OR3x1_ASAP7_75t_R register___U11702 ( .A(register__n350), .B(register__n7677), .C(register__n7676), .Y(register__n10975) );
  OA22x2_ASAP7_75t_R register___U11703 ( .A1(register__n420), .A2(register__n5732), .B1(register__n800), .B2(register__n11584), 
        .Y(register__n10978) );
  INVx1_ASAP7_75t_R register___U11704 ( .A(register__n5630), .Y(register__n7676) );
  OA222x2_ASAP7_75t_R register___U11705 ( .A1(register__n2002), .A2(register__n5246), .B1(register__n1997), .B2(
        net113158), .C1(register__net112580), .C2(register__n11587), .Y(register__n10976) );
  OA22x2_ASAP7_75t_R register___U11706 ( .A1(register__n66), .A2(register__n6233), .B1(register__n1691), .B2(register__n7246), 
        .Y(register__n10977) );
  BUFx4f_ASAP7_75t_R register___U11707 ( .A(register__net108114), .Y(register__net104596) );
  BUFx4f_ASAP7_75t_R register___U11708 ( .A(register__net122333), .Y(register__net104592) );
  BUFx6f_ASAP7_75t_R register___U11709 ( .A(register__n7681), .Y(register__n7680) );
  BUFx4f_ASAP7_75t_R register___U11710 ( .A(register__n5367), .Y(register__n7681) );
  BUFx6f_ASAP7_75t_R register___U11711 ( .A(register__n7683), .Y(register__n7682) );
  BUFx4f_ASAP7_75t_R register___U11712 ( .A(register__n6958), .Y(register__n7683) );
  BUFx4f_ASAP7_75t_R register___U11713 ( .A(register__net127327), .Y(register__net104579) );
  BUFx2_ASAP7_75t_R register___U11714 ( .A(register__n10598), .Y(register__n7688) );
  BUFx2_ASAP7_75t_R register___U11715 ( .A(register__n11348), .Y(register__n7689) );
  BUFx2_ASAP7_75t_R register___U11716 ( .A(register__n11203), .Y(register__n7690) );
  BUFx2_ASAP7_75t_R register___U11717 ( .A(register__n11179), .Y(register__n7691) );
  BUFx2_ASAP7_75t_R register___U11718 ( .A(register__n10575), .Y(register__n7692) );
  BUFx2_ASAP7_75t_R register___U11719 ( .A(register__C6422_net59856), .Y(register__net104283) );
  BUFx2_ASAP7_75t_R register___U11720 ( .A(register__n11128), .Y(register__n7693) );
  BUFx2_ASAP7_75t_R register___U11721 ( .A(register__n10741), .Y(register__n7694) );
  BUFx2_ASAP7_75t_R register___U11722 ( .A(register__n11663), .Y(register__n7695) );
  BUFx2_ASAP7_75t_R register___U11723 ( .A(register__n11061), .Y(register__n7696) );
  BUFx3_ASAP7_75t_R register___U11724 ( .A(register__n7699), .Y(register__n7698) );
  BUFx3_ASAP7_75t_R register___U11725 ( .A(register__n8033), .Y(register__n7702) );
  BUFx3_ASAP7_75t_R register___U11726 ( .A(register__n9702), .Y(register__n7703) );
  BUFx2_ASAP7_75t_R register___U11727 ( .A(register__n9702), .Y(register__n7704) );
  BUFx4f_ASAP7_75t_R register___U11728 ( .A(register__n9702), .Y(register__n7705) );
  BUFx3_ASAP7_75t_R register___U11729 ( .A(register__net98847), .Y(register__net104013) );
  BUFx3_ASAP7_75t_R register___U11730 ( .A(register__net98499), .Y(register__net104011) );
  BUFx12f_ASAP7_75t_R register___U11731 ( .A(register__n9781), .Y(register__n7707) );
  BUFx12f_ASAP7_75t_R register___U11732 ( .A(register__n9803), .Y(register__n7708) );
  BUFx3_ASAP7_75t_R register___U11733 ( .A(register__n9104), .Y(register__n7709) );
  BUFx12f_ASAP7_75t_R register___U11734 ( .A(register__net90258), .Y(register__net104001) );
  BUFx3_ASAP7_75t_R register___U11735 ( .A(register__net98215), .Y(register__net103999) );
  BUFx3_ASAP7_75t_R register___U11736 ( .A(register__n9134), .Y(register__n7710) );
  BUFx3_ASAP7_75t_R register___U11737 ( .A(register__n9138), .Y(register__n7711) );
  BUFx12f_ASAP7_75t_R register___U11738 ( .A(register__net88765), .Y(register__net103991) );
  BUFx3_ASAP7_75t_R register___U11739 ( .A(register__net94818), .Y(register__net103992) );
  BUFx12f_ASAP7_75t_R register___U11740 ( .A(register__net88761), .Y(register__net103987) );
  BUFx3_ASAP7_75t_R register___U11741 ( .A(register__net94810), .Y(register__net103988) );
  BUFx3_ASAP7_75t_R register___U11742 ( .A(register__net94776), .Y(register__net103985) );
  BUFx12f_ASAP7_75t_R register___U11743 ( .A(register__net88753), .Y(register__net103981) );
  BUFx3_ASAP7_75t_R register___U11744 ( .A(register__net94768), .Y(register__net103982) );
  BUFx3_ASAP7_75t_R register___U11745 ( .A(register__n8211), .Y(register__n7712) );
  BUFx2_ASAP7_75t_R register___U11746 ( .A(Reg_data[833]), .Y(register__n7713) );
  BUFx2_ASAP7_75t_R register___U11747 ( .A(Reg_data[832]), .Y(register__n7714) );
  BUFx2_ASAP7_75t_R register___U11748 ( .A(Reg_data[267]), .Y(register__net103947) );
  BUFx2_ASAP7_75t_R register___U11749 ( .A(Reg_data[271]), .Y(register__net103939) );
  BUFx6f_ASAP7_75t_R register___U11750 ( .A(register__net97169), .Y(register__net103940) );
  BUFx3_ASAP7_75t_R register___U11751 ( .A(register__net97169), .Y(register__net103941) );
  BUFx6f_ASAP7_75t_R register___U11752 ( .A(register__net97170), .Y(register__net97169) );
  BUFx4f_ASAP7_75t_R register___U11753 ( .A(register__net106310), .Y(register__net97170) );
  BUFx2_ASAP7_75t_R register___U11754 ( .A(Reg_data[275]), .Y(register__n7715) );
  BUFx2_ASAP7_75t_R register___U11755 ( .A(Reg_data[266]), .Y(register__net103924) );
  BUFx4f_ASAP7_75t_R register___U11756 ( .A(register__net103928), .Y(register__net103925) );
  BUFx6f_ASAP7_75t_R register___U11757 ( .A(register__net103927), .Y(register__net103926) );
  BUFx6f_ASAP7_75t_R register___U11758 ( .A(register__net97141), .Y(register__net103927) );
  BUFx3_ASAP7_75t_R register___U11759 ( .A(register__net97141), .Y(register__net103928) );
  BUFx6f_ASAP7_75t_R register___U11760 ( .A(register__net97142), .Y(register__net97141) );
  BUFx4f_ASAP7_75t_R register___U11761 ( .A(register__net106295), .Y(register__net97142) );
  BUFx2_ASAP7_75t_R register___U11762 ( .A(Reg_data[603]), .Y(register__n7716) );
  BUFx6f_ASAP7_75t_R register___U11763 ( .A(register__n8734), .Y(register__n7717) );
  BUFx3_ASAP7_75t_R register___U11764 ( .A(register__n8734), .Y(register__n7718) );
  BUFx6f_ASAP7_75t_R register___U11765 ( .A(register__n8735), .Y(register__n8734) );
  BUFx4f_ASAP7_75t_R register___U11766 ( .A(register__n6531), .Y(register__n8735) );
  BUFx2_ASAP7_75t_R register___U11767 ( .A(Reg_data[283]), .Y(register__n7719) );
  BUFx6f_ASAP7_75t_R register___U11768 ( .A(register__n8742), .Y(register__n7720) );
  BUFx3_ASAP7_75t_R register___U11769 ( .A(register__n8742), .Y(register__n7721) );
  BUFx6f_ASAP7_75t_R register___U11770 ( .A(register__n8743), .Y(register__n8742) );
  BUFx4f_ASAP7_75t_R register___U11771 ( .A(register__n6281), .Y(register__n8743) );
  BUFx2_ASAP7_75t_R register___U11772 ( .A(Reg_data[287]), .Y(register__n7722) );
  BUFx4f_ASAP7_75t_R register___U11773 ( .A(register__n7726), .Y(register__n7723) );
  BUFx6f_ASAP7_75t_R register___U11774 ( .A(register__n7725), .Y(register__n7724) );
  BUFx6f_ASAP7_75t_R register___U11775 ( .A(register__n9215), .Y(register__n7725) );
  BUFx3_ASAP7_75t_R register___U11776 ( .A(register__n9215), .Y(register__n7726) );
  INVx2_ASAP7_75t_R register___U11777 ( .A(register__n7724), .Y(register__n11129) );
  BUFx6f_ASAP7_75t_R register___U11778 ( .A(register__n9216), .Y(register__n9215) );
  BUFx4f_ASAP7_75t_R register___U11779 ( .A(register__n7379), .Y(register__n9216) );
  BUFx2_ASAP7_75t_R register___U11780 ( .A(Reg_data[351]), .Y(register__n7727) );
  BUFx2_ASAP7_75t_R register___U11781 ( .A(Reg_data[605]), .Y(register__net103891) );
  BUFx3_ASAP7_75t_R register___U11782 ( .A(register__net103752), .Y(register__net103751) );
  BUFx2_ASAP7_75t_R register___U11783 ( .A(Reg_data[966]), .Y(register__net103752) );
  BUFx3_ASAP7_75t_R register___U11784 ( .A(register__n7730), .Y(register__n7729) );
  BUFx2_ASAP7_75t_R register___U11785 ( .A(Reg_data[936]), .Y(register__n7730) );
  BUFx12f_ASAP7_75t_R register___U11786 ( .A(register__n9588), .Y(register__n7731) );
  BUFx12f_ASAP7_75t_R register___U11787 ( .A(register__n7731), .Y(register__n9587) );
  BUFx3_ASAP7_75t_R register___U11788 ( .A(register__n7733), .Y(register__n7732) );
  BUFx2_ASAP7_75t_R register___U11789 ( .A(Reg_data[899]), .Y(register__n7733) );
  BUFx3_ASAP7_75t_R register___U11790 ( .A(register__n7735), .Y(register__n7734) );
  BUFx2_ASAP7_75t_R register___U11791 ( .A(Reg_data[898]), .Y(register__n7735) );
  BUFx4f_ASAP7_75t_R register___U11792 ( .A(register__n6808), .Y(register__n7736) );
  BUFx2_ASAP7_75t_R register___U11793 ( .A(Reg_data[820]), .Y(register__n7737) );
  BUFx12f_ASAP7_75t_R register___U11794 ( .A(register__n9612), .Y(register__n7738) );
  BUFx12f_ASAP7_75t_R register___U11795 ( .A(register__n7738), .Y(register__n9611) );
  BUFx6f_ASAP7_75t_R register___U11796 ( .A(register__n7736), .Y(register__n9612) );
  BUFx3_ASAP7_75t_R register___U11797 ( .A(register__n7740), .Y(register__n7739) );
  BUFx2_ASAP7_75t_R register___U11798 ( .A(Reg_data[449]), .Y(register__n7740) );
  BUFx3_ASAP7_75t_R register___U11799 ( .A(register__net103721), .Y(register__net103720) );
  BUFx2_ASAP7_75t_R register___U11800 ( .A(Reg_data[389]), .Y(register__net103721) );
  BUFx3_ASAP7_75t_R register___U11801 ( .A(register__n7742), .Y(register__n7741) );
  BUFx2_ASAP7_75t_R register___U11802 ( .A(Reg_data[388]), .Y(register__n7742) );
  BUFx3_ASAP7_75t_R register___U11803 ( .A(register__n7744), .Y(register__n7743) );
  BUFx2_ASAP7_75t_R register___U11804 ( .A(Reg_data[338]), .Y(register__n7744) );
  BUFx3_ASAP7_75t_R register___U11805 ( .A(register__net103709), .Y(register__net103708) );
  BUFx2_ASAP7_75t_R register___U11806 ( .A(Reg_data[325]), .Y(register__net103709) );
  BUFx3_ASAP7_75t_R register___U11807 ( .A(register__n7746), .Y(register__n7745) );
  BUFx2_ASAP7_75t_R register___U11808 ( .A(Reg_data[320]), .Y(register__n7746) );
  BUFx3_ASAP7_75t_R register___U11809 ( .A(register__n7748), .Y(register__n7747) );
  BUFx2_ASAP7_75t_R register___U11810 ( .A(Reg_data[310]), .Y(register__n7748) );
  BUFx3_ASAP7_75t_R register___U11811 ( .A(register__n7750), .Y(register__n7749) );
  BUFx2_ASAP7_75t_R register___U11812 ( .A(Reg_data[309]), .Y(register__n7750) );
  BUFx3_ASAP7_75t_R register___U11813 ( .A(register__n7752), .Y(register__n7751) );
  BUFx2_ASAP7_75t_R register___U11814 ( .A(Reg_data[306]), .Y(register__n7752) );
  BUFx3_ASAP7_75t_R register___U11815 ( .A(register__n7754), .Y(register__n7753) );
  BUFx2_ASAP7_75t_R register___U11816 ( .A(Reg_data[304]), .Y(register__n7754) );
  BUFx3_ASAP7_75t_R register___U11817 ( .A(register__n7756), .Y(register__n7755) );
  BUFx2_ASAP7_75t_R register___U11818 ( .A(Reg_data[292]), .Y(register__n7756) );
  BUFx3_ASAP7_75t_R register___U11819 ( .A(register__n7758), .Y(register__n7757) );
  BUFx2_ASAP7_75t_R register___U11820 ( .A(Reg_data[290]), .Y(register__n7758) );
  BUFx3_ASAP7_75t_R register___U11821 ( .A(register__n7760), .Y(register__n7759) );
  BUFx2_ASAP7_75t_R register___U11822 ( .A(Reg_data[288]), .Y(register__n7760) );
  BUFx3_ASAP7_75t_R register___U11823 ( .A(register__n7762), .Y(register__n7761) );
  BUFx2_ASAP7_75t_R register___U11824 ( .A(Reg_data[277]), .Y(register__n7762) );
  BUFx3_ASAP7_75t_R register___U11825 ( .A(register__net103669), .Y(register__net103668) );
  BUFx2_ASAP7_75t_R register___U11826 ( .A(Reg_data[185]), .Y(register__net103669) );
  BUFx2_ASAP7_75t_R register___U11827 ( .A(Reg_data[180]), .Y(register__n7764) );
  BUFx3_ASAP7_75t_R register___U11828 ( .A(register__n7766), .Y(register__n7765) );
  BUFx2_ASAP7_75t_R register___U11829 ( .A(Reg_data[162]), .Y(register__n7766) );
  BUFx3_ASAP7_75t_R register___U11830 ( .A(register__n7768), .Y(register__n7767) );
  BUFx2_ASAP7_75t_R register___U11831 ( .A(Reg_data[65]), .Y(register__n7768) );
  BUFx3_ASAP7_75t_R register___U11832 ( .A(register__net103650), .Y(register__net103649) );
  BUFx2_ASAP7_75t_R register___U11833 ( .A(Reg_data[5]), .Y(register__net103650) );
  BUFx3_ASAP7_75t_R register___U11834 ( .A(register__n7770), .Y(register__n7769) );
  BUFx2_ASAP7_75t_R register___U11835 ( .A(Reg_data[246]), .Y(register__n7770) );
  BUFx3_ASAP7_75t_R register___U11836 ( .A(register__net103642), .Y(register__net103641) );
  BUFx2_ASAP7_75t_R register___U11837 ( .A(Reg_data[38]), .Y(register__net103642) );
  BUFx2_ASAP7_75t_R register___U11838 ( .A(Reg_data[232]), .Y(register__n7772) );
  BUFx3_ASAP7_75t_R register___U11839 ( .A(register__net103631), .Y(register__net103630) );
  BUFx2_ASAP7_75t_R register___U11840 ( .A(Reg_data[230]), .Y(register__net103631) );
  BUFx3_ASAP7_75t_R register___U11841 ( .A(register__n7774), .Y(register__n7773) );
  BUFx2_ASAP7_75t_R register___U11842 ( .A(Reg_data[228]), .Y(register__n7774) );
  BUFx3_ASAP7_75t_R register___U11843 ( .A(register__net103623), .Y(register__net103622) );
  BUFx2_ASAP7_75t_R register___U11844 ( .A(Reg_data[587]), .Y(register__net103623) );
  BUFx3_ASAP7_75t_R register___U11845 ( .A(register__n7776), .Y(register__n7775) );
  BUFx2_ASAP7_75t_R register___U11846 ( .A(Reg_data[45]), .Y(register__n7776) );
  BUFx3_ASAP7_75t_R register___U11847 ( .A(register__net103612), .Y(register__net103611) );
  BUFx2_ASAP7_75t_R register___U11848 ( .A(Reg_data[171]), .Y(register__net103612) );
  BUFx3_ASAP7_75t_R register___U11849 ( .A(register__n7778), .Y(register__n7777) );
  BUFx2_ASAP7_75t_R register___U11850 ( .A(Reg_data[590]), .Y(register__n7778) );
  BUFx12f_ASAP7_75t_R register___U11851 ( .A(register__n7780), .Y(register__n7779) );
  BUFx12f_ASAP7_75t_R register___U11852 ( .A(register__n9528), .Y(register__n7780) );
  BUFx3_ASAP7_75t_R register___U11853 ( .A(register__n7782), .Y(register__n7781) );
  BUFx2_ASAP7_75t_R register___U11854 ( .A(Reg_data[595]), .Y(register__n7782) );
  BUFx3_ASAP7_75t_R register___U11855 ( .A(register__n7784), .Y(register__n7783) );
  BUFx2_ASAP7_75t_R register___U11856 ( .A(Reg_data[237]), .Y(register__n7784) );
  BUFx3_ASAP7_75t_R register___U11857 ( .A(register__n7786), .Y(register__n7785) );
  BUFx2_ASAP7_75t_R register___U11858 ( .A(Reg_data[382]), .Y(register__n7786) );
  BUFx3_ASAP7_75t_R register___U11859 ( .A(register__n7788), .Y(register__n7787) );
  BUFx2_ASAP7_75t_R register___U11860 ( .A(Reg_data[295]), .Y(register__n7788) );
  BUFx12f_ASAP7_75t_R register___U11861 ( .A(register__n9763), .Y(register__n7789) );
  BUFx12f_ASAP7_75t_R register___U11862 ( .A(register__n7789), .Y(register__n9762) );
  BUFx3_ASAP7_75t_R register___U11863 ( .A(register__net103581), .Y(register__net103580) );
  BUFx2_ASAP7_75t_R register___U11864 ( .A(Reg_data[280]), .Y(register__net103581) );
  BUFx3_ASAP7_75t_R register___U11865 ( .A(register__n7791), .Y(register__n7790) );
  BUFx2_ASAP7_75t_R register___U11866 ( .A(Reg_data[334]), .Y(register__n7791) );
  BUFx3_ASAP7_75t_R register___U11867 ( .A(register__net103567), .Y(register__net103566) );
  BUFx2_ASAP7_75t_R register___U11868 ( .A(Reg_data[216]), .Y(register__net103567) );
  BUFx4f_ASAP7_75t_R register___U11869 ( .A(register__net89417), .Y(register__net103568) );
  BUFx2_ASAP7_75t_R register___U11870 ( .A(register__net89417), .Y(register__net103569) );
  BUFx3_ASAP7_75t_R register___U11871 ( .A(register__net103557), .Y(register__net103556) );
  BUFx2_ASAP7_75t_R register___U11872 ( .A(Reg_data[815]), .Y(register__net103557) );
  BUFx2_ASAP7_75t_R register___U11873 ( .A(register__net90533), .Y(register__net103558) );
  BUFx4f_ASAP7_75t_R register___U11874 ( .A(register__net90533), .Y(register__net103560) );
  BUFx3_ASAP7_75t_R register___U11875 ( .A(register__net103553), .Y(register__net103552) );
  BUFx2_ASAP7_75t_R register___U11876 ( .A(Reg_data[207]), .Y(register__net103553) );
  BUFx3_ASAP7_75t_R register___U11877 ( .A(register__n7793), .Y(register__n7792) );
  BUFx2_ASAP7_75t_R register___U11878 ( .A(Reg_data[19]), .Y(register__n7793) );
  BUFx3_ASAP7_75t_R register___U11879 ( .A(register__net103541), .Y(register__net103540) );
  BUFx2_ASAP7_75t_R register___U11880 ( .A(Reg_data[586]), .Y(register__net103541) );
  BUFx12f_ASAP7_75t_R register___U11881 ( .A(register__net103543), .Y(register__net103542) );
  BUFx12f_ASAP7_75t_R register___U11882 ( .A(register__net91220), .Y(register__net103543) );
  BUFx3_ASAP7_75t_R register___U11883 ( .A(register__n7795), .Y(register__n7794) );
  BUFx2_ASAP7_75t_R register___U11884 ( .A(Reg_data[435]), .Y(register__n7795) );
  BUFx3_ASAP7_75t_R register___U11885 ( .A(register__n7797), .Y(register__n7796) );
  BUFx2_ASAP7_75t_R register___U11886 ( .A(Reg_data[268]), .Y(register__n7797) );
  BUFx3_ASAP7_75t_R register___U11887 ( .A(register__n7799), .Y(register__n7798) );
  BUFx2_ASAP7_75t_R register___U11888 ( .A(Reg_data[935]), .Y(register__n7799) );
  BUFx3_ASAP7_75t_R register___U11889 ( .A(register__n9784), .Y(register__n7800) );
  BUFx6f_ASAP7_75t_R register___U11890 ( .A(register__n9784), .Y(register__n7801) );
  BUFx3_ASAP7_75t_R register___U11891 ( .A(register__n7803), .Y(register__n7802) );
  BUFx2_ASAP7_75t_R register___U11892 ( .A(Reg_data[636]), .Y(register__n7803) );
  BUFx3_ASAP7_75t_R register___U11893 ( .A(register__n7805), .Y(register__n7804) );
  BUFx2_ASAP7_75t_R register___U11894 ( .A(Reg_data[585]), .Y(register__n7805) );
  BUFx3_ASAP7_75t_R register___U11895 ( .A(register__n7807), .Y(register__n7806) );
  BUFx2_ASAP7_75t_R register___U11896 ( .A(Reg_data[302]), .Y(register__n7807) );
  BUFx3_ASAP7_75t_R register___U11897 ( .A(register__n9790), .Y(register__n7808) );
  BUFx2_ASAP7_75t_R register___U11898 ( .A(register__n9790), .Y(register__n7809) );
  BUFx4f_ASAP7_75t_R register___U11899 ( .A(register__n9790), .Y(register__n7810) );
  BUFx2_ASAP7_75t_R register___U11900 ( .A(Reg_data[174]), .Y(register__n7812) );
  BUFx3_ASAP7_75t_R register___U11901 ( .A(register__n7814), .Y(register__n7813) );
  BUFx2_ASAP7_75t_R register___U11902 ( .A(Reg_data[846]), .Y(register__n7814) );
  BUFx3_ASAP7_75t_R register___U11903 ( .A(register__n7816), .Y(register__n7815) );
  BUFx2_ASAP7_75t_R register___U11904 ( .A(Reg_data[92]), .Y(register__n7816) );
  BUFx3_ASAP7_75t_R register___U11905 ( .A(register__n7818), .Y(register__n7817) );
  BUFx2_ASAP7_75t_R register___U11906 ( .A(Reg_data[284]), .Y(register__n7818) );
  BUFx3_ASAP7_75t_R register___U11907 ( .A(register__n7820), .Y(register__n7819) );
  BUFx2_ASAP7_75t_R register___U11908 ( .A(Reg_data[467]), .Y(register__n7820) );
  BUFx4f_ASAP7_75t_R register___U11909 ( .A(register__n9818), .Y(register__n7821) );
  BUFx2_ASAP7_75t_R register___U11910 ( .A(register__n9818), .Y(register__n7822) );
  BUFx2_ASAP7_75t_R register___U11911 ( .A(register__n9818), .Y(register__n7823) );
  BUFx3_ASAP7_75t_R register___U11912 ( .A(register__n7825), .Y(register__n7824) );
  BUFx2_ASAP7_75t_R register___U11913 ( .A(Reg_data[339]), .Y(register__n7825) );
  BUFx3_ASAP7_75t_R register___U11914 ( .A(register__net103464), .Y(register__net103463) );
  BUFx2_ASAP7_75t_R register___U11915 ( .A(Reg_data[298]), .Y(register__net103464) );
  BUFx2_ASAP7_75t_R register___U11916 ( .A(register__net90405), .Y(register__net103466) );
  BUFx4f_ASAP7_75t_R register___U11917 ( .A(register__net90405), .Y(register__net103467) );
  BUFx3_ASAP7_75t_R register___U11918 ( .A(register__net103454), .Y(register__net103453) );
  BUFx2_ASAP7_75t_R register___U11919 ( .A(Reg_data[202]), .Y(register__net103454) );
  BUFx4f_ASAP7_75t_R register___U11920 ( .A(register__net89205), .Y(register__net103455) );
  BUFx2_ASAP7_75t_R register___U11921 ( .A(register__net89205), .Y(register__net103457) );
  BUFx3_ASAP7_75t_R register___U11922 ( .A(register__net103450), .Y(register__net103449) );
  BUFx2_ASAP7_75t_R register___U11923 ( .A(Reg_data[74]), .Y(register__net103450) );
  BUFx4f_ASAP7_75t_R register___U11924 ( .A(register__net106293), .Y(register__net103439) );
  BUFx12f_ASAP7_75t_R register___U11925 ( .A(register__net103442), .Y(register__net96598) );
  BUFx12f_ASAP7_75t_R register___U11926 ( .A(register__net96599), .Y(register__net103442) );
  BUFx6f_ASAP7_75t_R register___U11927 ( .A(register__net103439), .Y(register__net96599) );
  BUFx3_ASAP7_75t_R register___U11928 ( .A(register__n7827), .Y(register__n7826) );
  BUFx2_ASAP7_75t_R register___U11929 ( .A(Reg_data[183]), .Y(register__n7827) );
  BUFx12f_ASAP7_75t_R register___U11930 ( .A(register__n10254), .Y(register__n7828) );
  BUFx12f_ASAP7_75t_R register___U11931 ( .A(register__n7828), .Y(register__n10253) );
  BUFx3_ASAP7_75t_R register___U11932 ( .A(register__n7830), .Y(register__n7829) );
  BUFx2_ASAP7_75t_R register___U11933 ( .A(Reg_data[763]), .Y(register__n7830) );
  BUFx3_ASAP7_75t_R register___U11934 ( .A(register__n7832), .Y(register__n7831) );
  BUFx2_ASAP7_75t_R register___U11935 ( .A(Reg_data[311]), .Y(register__n7832) );
  BUFx3_ASAP7_75t_R register___U11936 ( .A(register__n7834), .Y(register__n7833) );
  BUFx2_ASAP7_75t_R register___U11937 ( .A(Reg_data[73]), .Y(register__n7834) );
  BUFx3_ASAP7_75t_R register___U11938 ( .A(register__n7836), .Y(register__n7835) );
  BUFx2_ASAP7_75t_R register___U11939 ( .A(Reg_data[329]), .Y(register__n7836) );
  BUFx3_ASAP7_75t_R register___U11940 ( .A(register__n7838), .Y(register__n7837) );
  BUFx2_ASAP7_75t_R register___U11941 ( .A(Reg_data[666]), .Y(register__n7838) );
  BUFx3_ASAP7_75t_R register___U11942 ( .A(register__n7840), .Y(register__n7839) );
  BUFx2_ASAP7_75t_R register___U11943 ( .A(Reg_data[159]), .Y(register__n7840) );
  BUFx3_ASAP7_75t_R register___U11944 ( .A(register__n10293), .Y(register__n7841) );
  BUFx2_ASAP7_75t_R register___U11945 ( .A(register__n10293), .Y(register__n7842) );
  BUFx4f_ASAP7_75t_R register___U11946 ( .A(register__n10293), .Y(register__n7843) );
  BUFx3_ASAP7_75t_R register___U11947 ( .A(register__n7845), .Y(register__n7844) );
  BUFx2_ASAP7_75t_R register___U11948 ( .A(Reg_data[799]), .Y(register__n7845) );
  BUFx4f_ASAP7_75t_R register___U11949 ( .A(register__n7848), .Y(register__n7846) );
  BUFx6f_ASAP7_75t_R register___U11950 ( .A(register__n7849), .Y(register__n7847) );
  BUFx3_ASAP7_75t_R register___U11951 ( .A(register__n9377), .Y(register__n7848) );
  BUFx6f_ASAP7_75t_R register___U11952 ( .A(register__n9377), .Y(register__n7849) );
  INVx1_ASAP7_75t_R register___U11953 ( .A(register__n7847), .Y(register__n11127) );
  BUFx3_ASAP7_75t_R register___U11954 ( .A(register__n7851), .Y(register__n7850) );
  BUFx2_ASAP7_75t_R register___U11955 ( .A(Reg_data[76]), .Y(register__n7851) );
  BUFx4f_ASAP7_75t_R register___U11956 ( .A(register__n5179), .Y(register__n7852) );
  BUFx2_ASAP7_75t_R register___U11957 ( .A(Reg_data[945]), .Y(register__n7853) );
  BUFx12f_ASAP7_75t_R register___U11958 ( .A(register__n8348), .Y(register__n8347) );
  BUFx6f_ASAP7_75t_R register___U11959 ( .A(register__n7852), .Y(register__n8348) );
  BUFx3_ASAP7_75t_R register___U11960 ( .A(register__n7855), .Y(register__n7854) );
  BUFx2_ASAP7_75t_R register___U11961 ( .A(Reg_data[177]), .Y(register__n7855) );
  BUFx12f_ASAP7_75t_R register___U11962 ( .A(register__n8804), .Y(register__n7856) );
  BUFx12f_ASAP7_75t_R register___U11963 ( .A(register__n7856), .Y(register__n8803) );
  BUFx3_ASAP7_75t_R register___U11964 ( .A(register__net103365), .Y(register__net103364) );
  BUFx2_ASAP7_75t_R register___U11965 ( .A(Reg_data[824]), .Y(register__net103365) );
  BUFx3_ASAP7_75t_R register___U11966 ( .A(register__n7858), .Y(register__n7857) );
  BUFx2_ASAP7_75t_R register___U11967 ( .A(Reg_data[27]), .Y(register__n7858) );
  BUFx3_ASAP7_75t_R register___U11968 ( .A(register__n7860), .Y(register__n7859) );
  BUFx2_ASAP7_75t_R register___U11969 ( .A(Reg_data[91]), .Y(register__n7860) );
  BUFx3_ASAP7_75t_R register___U11970 ( .A(register__net103353), .Y(register__net103352) );
  BUFx2_ASAP7_75t_R register___U11971 ( .A(Reg_data[573]), .Y(register__net103353) );
  BUFx3_ASAP7_75t_R register___U11972 ( .A(register__n7862), .Y(register__n7861) );
  BUFx2_ASAP7_75t_R register___U11973 ( .A(Reg_data[414]), .Y(register__n7862) );
  BUFx3_ASAP7_75t_R register___U11974 ( .A(register__n7864), .Y(register__n7863) );
  BUFx2_ASAP7_75t_R register___U11975 ( .A(Reg_data[430]), .Y(register__n7864) );
  BUFx12f_ASAP7_75t_R register___U11976 ( .A(register__n9908), .Y(register__n7865) );
  BUFx12f_ASAP7_75t_R register___U11977 ( .A(register__n7865), .Y(register__n9907) );
  BUFx4f_ASAP7_75t_R register___U11978 ( .A(register__n11548), .Y(register__n7866) );
  INVx2_ASAP7_75t_R register___U11979 ( .A(register__n8716), .Y(register__n11548) );
  BUFx6f_ASAP7_75t_R register___U11980 ( .A(register__n8717), .Y(register__n8716) );
  INVx2_ASAP7_75t_R register___U11981 ( .A(register__net97161), .Y(register__net103314) );
  BUFx4f_ASAP7_75t_R register___U11982 ( .A(register__C6422_net60277), .Y(register__net103310) );
  INVx2_ASAP7_75t_R register___U11983 ( .A(register__net106157), .Y(register__C6422_net60277) );
  BUFx6f_ASAP7_75t_R register___U11984 ( .A(register__net97118), .Y(register__net97117) );
  INVx2_ASAP7_75t_R register___U11985 ( .A(register__n9211), .Y(register__n11526) );
  BUFx6f_ASAP7_75t_R register___U11986 ( .A(register__n9212), .Y(register__n9211) );
  INVx2_ASAP7_75t_R register___U11987 ( .A(register__net99940), .Y(register__net103300) );
  BUFx6f_ASAP7_75t_R register___U11988 ( .A(register__net99941), .Y(register__net99940) );
  BUFx2_ASAP7_75t_R register___U11989 ( .A(register__C6423_net60748), .Y(register__net103295) );
  BUFx6f_ASAP7_75t_R register___U11990 ( .A(register__net97178), .Y(register__net97177) );
  BUFx3_ASAP7_75t_R register___U11991 ( .A(register__n10786), .Y(register__n7868) );
  INVx2_ASAP7_75t_R register___U11992 ( .A(register__n7396), .Y(register__n10786) );
  BUFx6f_ASAP7_75t_R register___U11993 ( .A(register__n8731), .Y(register__n8730) );
  BUFx4f_ASAP7_75t_R register___U11994 ( .A(register__n11161), .Y(register__n7869) );
  INVx2_ASAP7_75t_R register___U11995 ( .A(register__n8714), .Y(register__n11161) );
  BUFx6f_ASAP7_75t_R register___U11996 ( .A(register__n8715), .Y(register__n8714) );
  BUFx4f_ASAP7_75t_R register___U11997 ( .A(register__n10868), .Y(register__n7870) );
  INVx2_ASAP7_75t_R register___U11998 ( .A(register__n8708), .Y(register__n10868) );
  BUFx6f_ASAP7_75t_R register___U11999 ( .A(register__n8709), .Y(register__n8708) );
  OA22x2_ASAP7_75t_R register___U12000 ( .A1(register__n12173), .A2(register__n2220), .B1(register__n10218), .B2(register__n3478), 
        .Y(register__n12788) );
  INVx1_ASAP7_75t_R register___U12001 ( .A(register__n4531), .Y(register__n7871) );
  OA22x2_ASAP7_75t_R register___U12002 ( .A1(register__net64438), .A2(register__n4267), .B1(register__net90457), .B2(
        n5184), .Y(register__n12626) );
  INVx4_ASAP7_75t_R register___U12003 ( .A(register__net64474), .Y(register__net64438) );
  OA22x2_ASAP7_75t_R register___U12004 ( .A1(register__net62674), .A2(register__n399), .B1(register__n10327), .B2(register__n3415), .Y(register__n13285) );
  INVx1_ASAP7_75t_R register___U12005 ( .A(register__n6256), .Y(register__n7872) );
  OA22x2_ASAP7_75t_R register___U12006 ( .A1(register__n12292), .A2(register__n4267), .B1(register__n9824), .B2(register__n11901), 
        .Y(register__n12617) );
  INVx1_ASAP7_75t_R register___U12007 ( .A(register__n4884), .Y(register__n7873) );
  OA22x2_ASAP7_75t_R register___U12008 ( .A1(register__net62836), .A2(register__n2220), .B1(register__net89001), .B2(
        n4177), .Y(register__n12778) );
  CKINVDCx10_ASAP7_75t_R register___U12009 ( .A(register__n12350), .Y(register__n7874) );
  BUFx6f_ASAP7_75t_R register___U12010 ( .A(register__n7874), .Y(register__n12361) );
  BUFx6f_ASAP7_75t_R register___U12011 ( .A(register__n7874), .Y(register__n12357) );
  BUFx6f_ASAP7_75t_R register___U12012 ( .A(register__n7874), .Y(register__n12356) );
  BUFx6f_ASAP7_75t_R register___U12013 ( .A(register__n7874), .Y(register__n12363) );
  BUFx6f_ASAP7_75t_R register___U12014 ( .A(register__n7874), .Y(register__n12358) );
  INVx1_ASAP7_75t_R register___U12015 ( .A(register__n4284), .Y(register__n7875) );
  INVx1_ASAP7_75t_R register___U12016 ( .A(register__n5112), .Y(register__n7876) );
  AO22x2_ASAP7_75t_R register___U12017 ( .A1(register__n9278), .A2(register__net118097), .B1(register__n9931), .B2(
        net150890), .Y(register__n11537) );
  INVx1_ASAP7_75t_R register___U12018 ( .A(register__n3056), .Y(register__n7880) );
  INVx1_ASAP7_75t_R register___U12019 ( .A(register__n3232), .Y(register__n7883) );
  INVx1_ASAP7_75t_R register___U12020 ( .A(register__n3114), .Y(register__n7885) );
  INVx1_ASAP7_75t_R register___U12021 ( .A(register__n3116), .Y(register__n7886) );
  OA22x2_ASAP7_75t_R register___U12022 ( .A1(register__net63322), .A2(register__n399), .B1(register__n10128), .B2(
        n11741), .Y(register__n13293) );
  INVx1_ASAP7_75t_R register___U12023 ( .A(register__n6247), .Y(register__n7890) );
  OA22x2_ASAP7_75t_R register___U12024 ( .A1(register__net63238), .A2(register__n399), .B1(register__net89645), .B2(
        n8335), .Y(register__n13292) );
  OA22x2_ASAP7_75t_R register___U12025 ( .A1(register__n12406), .A2(register__n11900), .B1(register__n9732), .B2(register__n11820), .Y(register__n12610) );
  OA22x2_ASAP7_75t_R register___U12026 ( .A1(register__n3253), .A2(register__n11900), .B1(register__n9738), .B2(register__n6139), 
        .Y(register__n12624) );
  OA22x2_ASAP7_75t_R register___U12027 ( .A1(register__n12200), .A2(register__n109), .B1(register__n9361), .B2(register__n6301), 
        .Y(register__n12844) );
  INVx1_ASAP7_75t_R register___U12028 ( .A(register__n7122), .Y(register__n7891) );
  OA22x2_ASAP7_75t_R register___U12029 ( .A1(register__net64768), .A2(register__n2220), .B1(register__net90113), .B2(
        n11805), .Y(register__n12794) );
  INVx1_ASAP7_75t_R register___U12030 ( .A(register__n4501), .Y(register__n7893) );
  OA22x2_ASAP7_75t_R register___U12031 ( .A1(register__n3593), .A2(register__n2220), .B1(register__n9939), .B2(register__n3477), 
        .Y(register__n12798) );
  INVx1_ASAP7_75t_R register___U12032 ( .A(register__n4503), .Y(register__n7895) );
  OA22x2_ASAP7_75t_R register___U12033 ( .A1(register__n12372), .A2(register__n109), .B1(register__n9953), .B2(register__n3021), 
        .Y(register__n12839) );
  INVx1_ASAP7_75t_R register___U12034 ( .A(register__n7118), .Y(register__n7896) );
  OA22x2_ASAP7_75t_R register___U12035 ( .A1(register__n5351), .A2(register__n109), .B1(register__n9957), .B2(register__n3452), 
        .Y(register__n12841) );
  INVx1_ASAP7_75t_R register___U12036 ( .A(register__n5004), .Y(register__n7897) );
  OA22x2_ASAP7_75t_R register___U12037 ( .A1(register__net63162), .A2(register__n1092), .B1(register__net90853), .B2(
        n11760), .Y(register__n13067) );
  INVx1_ASAP7_75t_R register___U12038 ( .A(register__n4653), .Y(register__n7898) );
  OA22x2_ASAP7_75t_R register___U12039 ( .A1(register__n12368), .A2(register__n1120), .B1(register__n9668), .B2(register__n11756), 
        .Y(register__n13070) );
  OA22x2_ASAP7_75t_R register___U12040 ( .A1(register__n12023), .A2(register__n1616), .B1(register__n9676), .B2(register__n3572), 
        .Y(register__n13085) );
  OA22x2_ASAP7_75t_R register___U12041 ( .A1(register__n12254), .A2(register__n399), .B1(register__n10038), .B2(register__n3349), 
        .Y(register__n13298) );
  INVx1_ASAP7_75t_R register___U12042 ( .A(register__n5964), .Y(register__n7899) );
  OA22x2_ASAP7_75t_R register___U12043 ( .A1(register__n5074), .A2(register__n399), .B1(register__n10042), .B2(register__n3417), 
        .Y(register__n13302) );
  INVx1_ASAP7_75t_R register___U12044 ( .A(register__n5966), .Y(register__n7900) );
  OA22x2_ASAP7_75t_R register___U12045 ( .A1(register__n12204), .A2(register__n4267), .B1(register__n9710), .B2(register__n3152), 
        .Y(register__n12620) );
  OA22x2_ASAP7_75t_R register___U12046 ( .A1(register__n12062), .A2(register__n4267), .B1(register__n9712), .B2(register__n5047), 
        .Y(register__n12628) );
  INVx1_ASAP7_75t_R register___U12047 ( .A(register__n5761), .Y(register__n7901) );
  OA22x2_ASAP7_75t_R register___U12048 ( .A1(register__n946), .A2(register__n4267), .B1(register__n9716), .B2(register__n11904), 
        .Y(register__n12633) );
  OA22x2_ASAP7_75t_R register___U12049 ( .A1(register__n12119), .A2(register__n109), .B1(register__n10110), .B2(register__n3021), 
        .Y(register__n12848) );
  OA22x2_ASAP7_75t_R register___U12050 ( .A1(register__net64430), .A2(register__n109), .B1(register__net89461), .B2(
        n11803), .Y(register__n12850) );
  OA22x2_ASAP7_75t_R register___U12051 ( .A1(register__n12089), .A2(register__n2220), .B1(register__n10169), .B2(register__n3261), 
        .Y(register__n12791) );
  OA22x2_ASAP7_75t_R register___U12052 ( .A1(register__net62844), .A2(register__n3159), .B1(register__net90217), .B2(
        n1540), .Y(register__n12581) );
  OA22x2_ASAP7_75t_R register___U12053 ( .A1(register__net62816), .A2(register__n3119), .B1(register__net89445), .B2(
        n5342), .Y(register__n13287) );
  INVx1_ASAP7_75t_R register___U12054 ( .A(register__n6510), .Y(register__n7905) );
  OA22x2_ASAP7_75t_R register___U12055 ( .A1(register__net62842), .A2(register__n11900), .B1(register__net94801), .B2(
        n3327), .Y(register__n12608) );
  BUFx12f_ASAP7_75t_R register___U12056 ( .A(register__net102927), .Y(register__net102924) );
  BUFx6f_ASAP7_75t_R register___U12057 ( .A(register__net102923), .Y(register__net64892) );
  BUFx6f_ASAP7_75t_R register___U12058 ( .A(register__n5185), .Y(register__n12239) );
  BUFx6f_ASAP7_75t_R register___U12059 ( .A(register__net64056), .Y(register__net64028) );
  BUFx12f_ASAP7_75t_R register___U12060 ( .A(register__n3727), .Y(register__n7907) );
  BUFx6f_ASAP7_75t_R register___U12061 ( .A(register__n12475), .Y(register__n12479) );
  INVx1_ASAP7_75t_R register___U12062 ( .A(register__n5021), .Y(register__n7910) );
  INVx1_ASAP7_75t_R register___U12063 ( .A(register__n5022), .Y(register__n7911) );
  INVx1_ASAP7_75t_R register___U12064 ( .A(register__n10947), .Y(register__n7912) );
  INVx1_ASAP7_75t_R register___U12065 ( .A(register__n4797), .Y(register__n7913) );
  INVx1_ASAP7_75t_R register___U12066 ( .A(register__n4799), .Y(register__n7914) );
  INVx1_ASAP7_75t_R register___U12067 ( .A(register__n5290), .Y(register__n7916) );
  INVx1_ASAP7_75t_R register___U12068 ( .A(register__n5292), .Y(register__n7917) );
  INVx1_ASAP7_75t_R register___U12069 ( .A(register__n5294), .Y(register__n7918) );
  INVx1_ASAP7_75t_R register___U12070 ( .A(register__n4570), .Y(register__n7919) );
  AND4x1_ASAP7_75t_R register___U12071 ( .A(register__n7920), .B(register__n1571), .C(register__n7922), .D(register__n4572), .Y(
        n11639) );
  AO22x1_ASAP7_75t_R register___U12072 ( .A1(register__n9599), .A2(register__n128), .B1(register__n10022), .B2(register__n1450), 
        .Y(register__n11439) );
  INVx1_ASAP7_75t_R register___U12073 ( .A(register__n5072), .Y(register__n7922) );
  INVx1_ASAP7_75t_R register___U12074 ( .A(register__n4306), .Y(register__n7923) );
  INVx1_ASAP7_75t_R register___U12075 ( .A(register__n4684), .Y(register__n7926) );
  INVx1_ASAP7_75t_R register___U12076 ( .A(register__n4686), .Y(register__n7927) );
  INVx1_ASAP7_75t_R register___U12077 ( .A(register__n5589), .Y(register__n7929) );
  INVx1_ASAP7_75t_R register___U12078 ( .A(register__n4701), .Y(register__n7930) );
  INVx1_ASAP7_75t_R register___U12079 ( .A(register__n11355), .Y(register__n7931) );
  INVx1_ASAP7_75t_R register___U12080 ( .A(register__n4612), .Y(register__n7932) );
  INVx1_ASAP7_75t_R register___U12081 ( .A(register__n4614), .Y(register__n7933) );
  INVx1_ASAP7_75t_R register___U12082 ( .A(register__n4723), .Y(register__n7934) );
  INVx1_ASAP7_75t_R register___U12083 ( .A(register__n3064), .Y(register__n7937) );
  BUFx2_ASAP7_75t_R register___U12084 ( .A(register__n10781), .Y(register__n7943) );
  INVx1_ASAP7_75t_R register___U12085 ( .A(register__n3630), .Y(register__n7944) );
  INVx1_ASAP7_75t_R register___U12086 ( .A(register__n3635), .Y(register__n7946) );
  INVx1_ASAP7_75t_R register___U12087 ( .A(register__n5623), .Y(register__n7947) );
  INVx1_ASAP7_75t_R register___U12088 ( .A(register__n5625), .Y(register__n7948) );
  AND4x1_ASAP7_75t_R register___U12089 ( .A(register__n1457), .B(register__n7947), .C(register__net100454), .D(register__n5627), 
        .Y(register__n11474) );
  OA22x2_ASAP7_75t_R register___U12090 ( .A1(register__n12315), .A2(register__n1092), .B1(register__n9672), .B2(register__n3822), 
        .Y(register__n13072) );
  OA22x2_ASAP7_75t_R register___U12091 ( .A1(register__net120805), .A2(register__n1120), .B1(register__net90833), .B2(
        n417), .Y(register__n13083) );
  OA22x2_ASAP7_75t_R register___U12092 ( .A1(register__n12175), .A2(register__n1092), .B1(register__n9758), .B2(register__n11759), 
        .Y(register__n13077) );
  OA22x2_ASAP7_75t_R register___U12093 ( .A1(register__net63004), .A2(register__n2220), .B1(register__n8793), .B2(register__n1462), .Y(register__n12780) );
  OA22x2_ASAP7_75t_R register___U12094 ( .A1(register__n12020), .A2(register__n11859), .B1(register__n10046), .B2(register__n3651), .Y(register__n13304) );
  OA22x2_ASAP7_75t_R register___U12095 ( .A1(register__n12455), .A2(register__n1755), .B1(register__n9788), .B2(register__n3821), 
        .Y(register__n13117) );
  INVx1_ASAP7_75t_R register___U12096 ( .A(register__n7356), .Y(register__n7951) );
  OA22x2_ASAP7_75t_R register___U12097 ( .A1(register__n3304), .A2(register__n1092), .B1(register__n10436), .B2(register__n3510), 
        .Y(register__n13066) );
  INVx1_ASAP7_75t_R register___U12098 ( .A(register__n13066), .Y(register__n7952) );
  OA22x2_ASAP7_75t_R register___U12099 ( .A1(register__n12424), .A2(register__n1755), .B1(register__n9349), .B2(register__n3821), 
        .Y(register__n13119) );
  OA22x2_ASAP7_75t_R register___U12100 ( .A1(register__n3319), .A2(register__n576), .B1(register__n5836), .B2(register__n585), 
        .Y(register__n13211) );
  INVx1_ASAP7_75t_R register___U12101 ( .A(register__n4529), .Y(register__n7953) );
  OA22x2_ASAP7_75t_R register___U12102 ( .A1(register__n420), .A2(register__n8360), .B1(register__n800), .B2(register__n11327), 
        .Y(register__n10660) );
  OA22x2_ASAP7_75t_R register___U12103 ( .A1(register__net107674), .A2(register__n7247), .B1(register__n1691), .B2(
        n6984), .Y(register__n10659) );
  INVx1_ASAP7_75t_R register___U12104 ( .A(register__n4930), .Y(register__n7957) );
  OA222x2_ASAP7_75t_R register___U12105 ( .A1(register__n2081), .A2(register__n5549), .B1(register__n817), .B2(register__n6470), 
        .C1(register__net112580), .C2(register__n9156), .Y(register__n10658) );
  OR3x1_ASAP7_75t_R register___U12106 ( .A(register__n7961), .B(register__n293), .C(register__n7960), .Y(register__n11563) );
  INVx1_ASAP7_75t_R register___U12107 ( .A(register__n5315), .Y(register__n7959) );
  OA22x2_ASAP7_75t_R register___U12108 ( .A1(register__net131654), .A2(register__n6227), .B1(register__net130175), .B2(
        n6776), .Y(register__n11565) );
  INVx1_ASAP7_75t_R register___U12109 ( .A(register__n5316), .Y(register__n7960) );
  OA22x2_ASAP7_75t_R register___U12110 ( .A1(register__n713), .A2(register__n7340), .B1(register__net149937), .B2(
        n10957), .Y(register__n11564) );
  INVx1_ASAP7_75t_R register___U12111 ( .A(register__n5317), .Y(register__n7961) );
  OR3x1_ASAP7_75t_R register___U12112 ( .A(register__n5998), .B(register__n7964), .C(register__n7962), .Y(register__n11241) );
  OA22x2_ASAP7_75t_R register___U12113 ( .A1(register__net131654), .A2(register__n11245), .B1(register__net130175), 
        .B2(register__n6985), .Y(register__n11244) );
  INVx1_ASAP7_75t_R register___U12114 ( .A(register__n5996), .Y(register__n7962) );
  OA222x2_ASAP7_75t_R register___U12115 ( .A1(register__n1987), .A2(register__n10621), .B1(register__n1995), .B2(
        net112155), .C1(register__n1800), .C2(register__n6207), .Y(register__n11242) );
  OA22x2_ASAP7_75t_R register___U12116 ( .A1(register__n714), .A2(register__n7586), .B1(register__net149937), .B2(register__n7243), .Y(register__n11243) );
  OR3x1_ASAP7_75t_R register___U12117 ( .A(register__n4927), .B(register__n7966), .C(register__n7965), .Y(register__n10819) );
  INVx1_ASAP7_75t_R register___U12118 ( .A(register__n4923), .Y(register__n7965) );
  OA22x2_ASAP7_75t_R register___U12119 ( .A1(register__net107674), .A2(register__n11435), .B1(register__n1691), .B2(
        n8216), .Y(register__n10821) );
  INVx1_ASAP7_75t_R register___U12120 ( .A(register__n4925), .Y(register__n7966) );
  OA222x2_ASAP7_75t_R register___U12121 ( .A1(register__n1978), .A2(register__n6215), .B1(register__n817), .B2(register__n5724), 
        .C1(register__net112578), .C2(register__n11437), .Y(register__n10820) );
  INVx1_ASAP7_75t_R register___U12122 ( .A(register__n10820), .Y(register__n7967) );
  OA22x2_ASAP7_75t_R register___U12123 ( .A1(register__n420), .A2(register__n10760), .B1(register__n802), .B2(register__n6773), 
        .Y(register__n10759) );
  OA22x2_ASAP7_75t_R register___U12124 ( .A1(register__net107674), .A2(register__n8009), .B1(register__n1691), .B2(
        n7343), .Y(register__n10758) );
  OR3x1_ASAP7_75t_R register___U12125 ( .A(register__n5150), .B(register__n7969), .C(register__n7968), .Y(register__n11300) );
  OA22x2_ASAP7_75t_R register___U12126 ( .A1(register__net131654), .A2(register__n6482), .B1(register__net130175), .B2(
        n8362), .Y(register__n11303) );
  INVx1_ASAP7_75t_R register___U12127 ( .A(register__n5149), .Y(register__n7968) );
  OA22x2_ASAP7_75t_R register___U12128 ( .A1(register__n710), .A2(register__n9148), .B1(register__n353), .B2(register__n7245), 
        .Y(register__n11302) );
  OR3x1_ASAP7_75t_R register___U12129 ( .A(register__n6020), .B(register__n7971), .C(register__n7970), .Y(register__n11580) );
  OA22x2_ASAP7_75t_R register___U12130 ( .A1(register__net131654), .A2(register__n6774), .B1(register__net130175), .B2(
        n5733), .Y(register__n11582) );
  INVx1_ASAP7_75t_R register___U12131 ( .A(register__n6014), .Y(register__n7970) );
  OA22x2_ASAP7_75t_R register___U12132 ( .A1(register__n713), .A2(register__n6233), .B1(register__net149939), .B2(register__n7246), .Y(register__n11581) );
  INVx1_ASAP7_75t_R register___U12133 ( .A(register__n6016), .Y(register__n7971) );
  OR3x1_ASAP7_75t_R register___U12134 ( .A(register__n126), .B(register__n7975), .C(register__n7974), .Y(register__n10997) );
  OA22x2_ASAP7_75t_R register___U12135 ( .A1(register__n419), .A2(register__net113240), .B1(register__n800), .B2(
        net98142), .Y(register__n11000) );
  INVx1_ASAP7_75t_R register___U12136 ( .A(register__n5130), .Y(register__n7974) );
  OA22x2_ASAP7_75t_R register___U12137 ( .A1(register__net107674), .A2(register__net105496), .B1(register__n1691), .B2(
        net107815), .Y(register__n10999) );
  INVx1_ASAP7_75t_R register___U12138 ( .A(register__n5132), .Y(register__n7975) );
  OA222x2_ASAP7_75t_R register___U12139 ( .A1(register__n1978), .A2(register__C6423_net61141), .B1(register__n1997), 
        .B2(register__net117114), .C1(register__net112580), .C2(register__net109880), .Y(register__n10998) );
  OR3x1_ASAP7_75t_R register___U12140 ( .A(register__n558), .B(register__n7978), .C(register__n7977), .Y(register__n10841) );
  OA22x2_ASAP7_75t_R register___U12141 ( .A1(register__n420), .A2(register__n11454), .B1(register__n800), .B2(register__n11455), 
        .Y(register__n10844) );
  OA222x2_ASAP7_75t_R register___U12142 ( .A1(register__n2002), .A2(register__n6221), .B1(register__n1997), .B2(register__n10847), 
        .C1(register__net112580), .C2(register__n7575), .Y(register__n10842) );
  OA22x2_ASAP7_75t_R register___U12143 ( .A1(register__net107674), .A2(register__n6780), .B1(register__n1691), .B2(
        n7242), .Y(register__n10843) );
  INVx1_ASAP7_75t_R register___U12144 ( .A(register__n5147), .Y(register__n7978) );
  OR3x1_ASAP7_75t_R register___U12145 ( .A(register__n5827), .B(register__n7980), .C(register__n7979), .Y(register__n11618) );
  OA22x2_ASAP7_75t_R register___U12146 ( .A1(register__n2013), .A2(register__n6232), .B1(register__net130175), .B2(
        n9159), .Y(register__n11621) );
  INVx1_ASAP7_75t_R register___U12147 ( .A(register__n11621), .Y(register__n7979) );
  OA22x2_ASAP7_75t_R register___U12148 ( .A1(register__n710), .A2(register__register__n7107), .B1(register__net149934), .B2(register__n6489), .Y(register__n11620) );
  INVx1_ASAP7_75t_R register___U12149 ( .A(register__n5824), .Y(register__n7980) );
  INVx1_ASAP7_75t_R register___U12150 ( .A(register__n5826), .Y(register__n7981) );
  BUFx6f_ASAP7_75t_R register___U12151 ( .A(register__n7989), .Y(register__n7988) );
  BUFx4f_ASAP7_75t_R register___U12152 ( .A(register__n7432), .Y(register__n7989) );
  BUFx6f_ASAP7_75t_R register___U12153 ( .A(register__n7991), .Y(register__n7990) );
  BUFx4f_ASAP7_75t_R register___U12154 ( .A(register__n7445), .Y(register__n7991) );
  BUFx6f_ASAP7_75t_R register___U12155 ( .A(register__n7993), .Y(register__n7992) );
  BUFx4f_ASAP7_75t_R register___U12156 ( .A(register__n5895), .Y(register__n7993) );
  BUFx6f_ASAP7_75t_R register___U12157 ( .A(register__n7995), .Y(register__n7994) );
  BUFx4f_ASAP7_75t_R register___U12158 ( .A(register__n6328), .Y(register__n7995) );
  BUFx6f_ASAP7_75t_R register___U12159 ( .A(register__n7998), .Y(register__n7997) );
  BUFx4f_ASAP7_75t_R register___U12160 ( .A(register__n7505), .Y(register__n7998) );
  BUFx6f_ASAP7_75t_R register___U12161 ( .A(register__n8000), .Y(register__n7999) );
  BUFx4f_ASAP7_75t_R register___U12162 ( .A(register__n6951), .Y(register__n8000) );
  BUFx2_ASAP7_75t_R register___U12163 ( .A(register__n11326), .Y(register__n8001) );
  BUFx2_ASAP7_75t_R register___U12164 ( .A(register__C6423_net60617), .Y(register__net101833) );
  BUFx2_ASAP7_75t_R register___U12165 ( .A(register__n11201), .Y(register__n8002) );
  BUFx2_ASAP7_75t_R register___U12166 ( .A(register__n10595), .Y(register__n8003) );
  BUFx2_ASAP7_75t_R register___U12167 ( .A(register__n11394), .Y(register__n8004) );
  BUFx2_ASAP7_75t_R register___U12168 ( .A(register__n11103), .Y(register__n8005) );
  BUFx2_ASAP7_75t_R register___U12169 ( .A(register__n11454), .Y(register__n8006) );
  BUFx2_ASAP7_75t_R register___U12170 ( .A(register__n11062), .Y(register__n8007) );
  BUFx2_ASAP7_75t_R register___U12171 ( .A(register__n11686), .Y(register__n8008) );
  BUFx2_ASAP7_75t_R register___U12172 ( .A(register__n10762), .Y(register__n8009) );
  BUFx3_ASAP7_75t_R register___U12173 ( .A(register__n8011), .Y(register__n8010) );
  BUFx2_ASAP7_75t_R register___U12174 ( .A(register__n11054), .Y(register__n8011) );
  INVx6_ASAP7_75t_R register___U12175 ( .A(register__net63190), .Y(register__net63158) );
  BUFx12f_ASAP7_75t_R register___U12176 ( .A(register__net145202), .Y(register__net63190) );
  INVx1_ASAP7_75t_R register___U12177 ( .A(register__n11268), .Y(register__n8013) );
  BUFx6f_ASAP7_75t_R register___U12178 ( .A(register__n8015), .Y(register__n8014) );
  BUFx4f_ASAP7_75t_R register___U12179 ( .A(register__n10956), .Y(register__n8015) );
  BUFx12f_ASAP7_75t_R register___U12180 ( .A(register__net89846), .Y(register__net101570) );
  BUFx3_ASAP7_75t_R register___U12181 ( .A(register__net95351), .Y(register__net101568) );
  BUFx3_ASAP7_75t_R register___U12182 ( .A(register__n8967), .Y(register__n8016) );
  BUFx3_ASAP7_75t_R register___U12183 ( .A(register__net95274), .Y(register__net101564) );
  BUFx3_ASAP7_75t_R register___U12184 ( .A(register__n8990), .Y(register__n8017) );
  BUFx3_ASAP7_75t_R register___U12185 ( .A(register__n9003), .Y(register__n8019) );
  BUFx3_ASAP7_75t_R register___U12186 ( .A(register__n9015), .Y(register__n8020) );
  BUFx3_ASAP7_75t_R register___U12187 ( .A(register__n8374), .Y(register__n8021) );
  BUFx3_ASAP7_75t_R register___U12188 ( .A(register__n8476), .Y(register__n8022) );
  BUFx3_ASAP7_75t_R register___U12189 ( .A(register__n8496), .Y(register__n8023) );
  BUFx3_ASAP7_75t_R register___U12190 ( .A(register__n9067), .Y(register__n8024) );
  BUFx12f_ASAP7_75t_R register___U12191 ( .A(register__n10236), .Y(register__n8025) );
  BUFx12f_ASAP7_75t_R register___U12192 ( .A(register__n10304), .Y(register__n8026) );
  INVx2_ASAP7_75t_R register___U12193 ( .A(register__n8724), .Y(register__n10980) );
  BUFx6f_ASAP7_75t_R register___U12194 ( .A(register__n8725), .Y(register__n8724) );
  BUFx2_ASAP7_75t_R register___U12195 ( .A(Reg_data[584]), .Y(register__n8027) );
  BUFx2_ASAP7_75t_R register___U12196 ( .A(Reg_data[581]), .Y(register__net101470) );
  BUFx2_ASAP7_75t_R register___U12197 ( .A(Reg_data[118]), .Y(register__n8028) );
  BUFx3_ASAP7_75t_R register___U12198 ( .A(register__n10032), .Y(register__n8029) );
  BUFx2_ASAP7_75t_R register___U12199 ( .A(register__n10032), .Y(register__n8030) );
  BUFx4f_ASAP7_75t_R register___U12200 ( .A(register__n10032), .Y(register__n8031) );
  BUFx6f_ASAP7_75t_R register___U12201 ( .A(register__n10033), .Y(register__n10032) );
  BUFx4f_ASAP7_75t_R register___U12202 ( .A(register__n7371), .Y(register__n10033) );
  BUFx2_ASAP7_75t_R register___U12203 ( .A(Reg_data[114]), .Y(register__n8032) );
  BUFx6f_ASAP7_75t_R register___U12204 ( .A(register__n10039), .Y(register__n10038) );
  BUFx4f_ASAP7_75t_R register___U12205 ( .A(register__n7372), .Y(register__n10039) );
  BUFx2_ASAP7_75t_R register___U12206 ( .A(Reg_data[112]), .Y(register__n8033) );
  BUFx6f_ASAP7_75t_R register___U12207 ( .A(register__n10041), .Y(register__n10040) );
  BUFx4f_ASAP7_75t_R register___U12208 ( .A(register__n7702), .Y(register__n10041) );
  BUFx2_ASAP7_75t_R register___U12209 ( .A(Reg_data[102]), .Y(register__net101448) );
  BUFx4f_ASAP7_75t_R register___U12210 ( .A(register__net106320), .Y(register__net89817) );
  BUFx2_ASAP7_75t_R register___U12211 ( .A(Reg_data[98]), .Y(register__n8034) );
  BUFx6f_ASAP7_75t_R register___U12212 ( .A(register__n10049), .Y(register__n10048) );
  BUFx4f_ASAP7_75t_R register___U12213 ( .A(register__n7373), .Y(register__n10049) );
  INVx1_ASAP7_75t_R register___U12214 ( .A(register__n11091), .Y(register__n8035) );
  INVx1_ASAP7_75t_R register___U12215 ( .A(register__n4993), .Y(register__n8036) );
  BUFx12f_ASAP7_75t_R register___U12216 ( .A(register__net144157), .Y(register__net64724) );
  BUFx12f_ASAP7_75t_R register___U12217 ( .A(register__net136275), .Y(register__net64702) );
  BUFx3_ASAP7_75t_R register___U12218 ( .A(register__net101358), .Y(register__net101357) );
  BUFx2_ASAP7_75t_R register___U12219 ( .A(Reg_data[934]), .Y(register__net101358) );
  BUFx3_ASAP7_75t_R register___U12220 ( .A(register__net101354), .Y(register__net101353) );
  BUFx2_ASAP7_75t_R register___U12221 ( .A(Reg_data[678]), .Y(register__net101354) );
  BUFx3_ASAP7_75t_R register___U12222 ( .A(register__n8039), .Y(register__n8038) );
  BUFx2_ASAP7_75t_R register___U12223 ( .A(Reg_data[674]), .Y(register__n8039) );
  BUFx3_ASAP7_75t_R register___U12224 ( .A(register__n8041), .Y(register__n8040) );
  BUFx2_ASAP7_75t_R register___U12225 ( .A(Reg_data[628]), .Y(register__n8041) );
  BUFx3_ASAP7_75t_R register___U12226 ( .A(register__n8043), .Y(register__n8042) );
  BUFx2_ASAP7_75t_R register___U12227 ( .A(Reg_data[626]), .Y(register__n8043) );
  BUFx3_ASAP7_75t_R register___U12228 ( .A(register__n8045), .Y(register__n8044) );
  BUFx2_ASAP7_75t_R register___U12229 ( .A(Reg_data[598]), .Y(register__n8045) );
  BUFx3_ASAP7_75t_R register___U12230 ( .A(register__n8047), .Y(register__n8046) );
  BUFx2_ASAP7_75t_R register___U12231 ( .A(Reg_data[578]), .Y(register__n8047) );
  BUFx3_ASAP7_75t_R register___U12232 ( .A(register__n8049), .Y(register__n8048) );
  BUFx2_ASAP7_75t_R register___U12233 ( .A(Reg_data[402]), .Y(register__n8049) );
  BUFx3_ASAP7_75t_R register___U12234 ( .A(register__net101326), .Y(register__net101325) );
  BUFx2_ASAP7_75t_R register___U12235 ( .A(Reg_data[377]), .Y(register__net101326) );
  BUFx3_ASAP7_75t_R register___U12236 ( .A(register__n8051), .Y(register__n8050) );
  BUFx2_ASAP7_75t_R register___U12237 ( .A(Reg_data[374]), .Y(register__n8051) );
  BUFx3_ASAP7_75t_R register___U12238 ( .A(register__n8053), .Y(register__n8052) );
  BUFx2_ASAP7_75t_R register___U12239 ( .A(Reg_data[368]), .Y(register__n8053) );
  BUFx3_ASAP7_75t_R register___U12240 ( .A(register__net101314), .Y(register__net101313) );
  BUFx2_ASAP7_75t_R register___U12241 ( .A(Reg_data[358]), .Y(register__net101314) );
  BUFx3_ASAP7_75t_R register___U12242 ( .A(register__n8055), .Y(register__n8054) );
  BUFx2_ASAP7_75t_R register___U12243 ( .A(Reg_data[336]), .Y(register__n8055) );
  BUFx3_ASAP7_75t_R register___U12244 ( .A(register__net101306), .Y(register__net101305) );
  BUFx2_ASAP7_75t_R register___U12245 ( .A(Reg_data[326]), .Y(register__net101306) );
  BUFx3_ASAP7_75t_R register___U12246 ( .A(register__n8057), .Y(register__n8056) );
  BUFx2_ASAP7_75t_R register___U12247 ( .A(Reg_data[321]), .Y(register__n8057) );
  BUFx3_ASAP7_75t_R register___U12248 ( .A(register__n8059), .Y(register__n8058) );
  BUFx2_ASAP7_75t_R register___U12249 ( .A(Reg_data[278]), .Y(register__n8059) );
  BUFx3_ASAP7_75t_R register___U12250 ( .A(register__n8061), .Y(register__n8060) );
  BUFx2_ASAP7_75t_R register___U12251 ( .A(Reg_data[258]), .Y(register__n8061) );
  BUFx3_ASAP7_75t_R register___U12252 ( .A(register__n8063), .Y(register__n8062) );
  BUFx2_ASAP7_75t_R register___U12253 ( .A(Reg_data[181]), .Y(register__n8063) );
  BUFx3_ASAP7_75t_R register___U12254 ( .A(register__n8065), .Y(register__n8064) );
  BUFx2_ASAP7_75t_R register___U12255 ( .A(Reg_data[164]), .Y(register__n8065) );
  BUFx3_ASAP7_75t_R register___U12256 ( .A(register__n8067), .Y(register__n8066) );
  BUFx2_ASAP7_75t_R register___U12257 ( .A(Reg_data[161]), .Y(register__n8067) );
  BUFx3_ASAP7_75t_R register___U12258 ( .A(register__n8069), .Y(register__n8068) );
  BUFx2_ASAP7_75t_R register___U12259 ( .A(Reg_data[149]), .Y(register__n8069) );
  BUFx3_ASAP7_75t_R register___U12260 ( .A(register__net101274), .Y(register__net101273) );
  BUFx2_ASAP7_75t_R register___U12261 ( .A(Reg_data[134]), .Y(register__net101274) );
  BUFx3_ASAP7_75t_R register___U12262 ( .A(register__n8071), .Y(register__n8070) );
  BUFx2_ASAP7_75t_R register___U12263 ( .A(Reg_data[104]), .Y(register__n8071) );
  BUFx3_ASAP7_75t_R register___U12264 ( .A(register__n8073), .Y(register__n8072) );
  BUFx2_ASAP7_75t_R register___U12265 ( .A(Reg_data[16]), .Y(register__n8073) );
  BUFx3_ASAP7_75t_R register___U12266 ( .A(register__n8075), .Y(register__n8074) );
  BUFx2_ASAP7_75t_R register___U12267 ( .A(Reg_data[1]), .Y(register__n8075) );
  BUFx3_ASAP7_75t_R register___U12268 ( .A(register__n8077), .Y(register__n8076) );
  BUFx2_ASAP7_75t_R register___U12269 ( .A(Reg_data[192]), .Y(register__n8077) );
  BUFx3_ASAP7_75t_R register___U12270 ( .A(register__n8079), .Y(register__n8078) );
  BUFx2_ASAP7_75t_R register___U12271 ( .A(Reg_data[32]), .Y(register__n8079) );
  BUFx3_ASAP7_75t_R register___U12272 ( .A(register__n8081), .Y(register__n8080) );
  BUFx2_ASAP7_75t_R register___U12273 ( .A(Reg_data[36]), .Y(register__n8081) );
  BUFx4f_ASAP7_75t_R register___U12274 ( .A(register__n10082), .Y(register__n8082) );
  BUFx2_ASAP7_75t_R register___U12275 ( .A(register__n10082), .Y(register__n8083) );
  BUFx2_ASAP7_75t_R register___U12276 ( .A(register__n10082), .Y(register__n8084) );
  BUFx3_ASAP7_75t_R register___U12277 ( .A(register__n8086), .Y(register__n8085) );
  BUFx2_ASAP7_75t_R register___U12278 ( .A(Reg_data[242]), .Y(register__n8086) );
  BUFx2_ASAP7_75t_R register___U12279 ( .A(Reg_data[48]), .Y(register__n8088) );
  BUFx4f_ASAP7_75t_R register___U12280 ( .A(register__n6524), .Y(register__n8089) );
  BUFx2_ASAP7_75t_R register___U12281 ( .A(Reg_data[807]), .Y(register__n8090) );
  BUFx12f_ASAP7_75t_R register___U12282 ( .A(register__n9721), .Y(register__n8091) );
  BUFx12f_ASAP7_75t_R register___U12283 ( .A(register__n8091), .Y(register__n9720) );
  BUFx6f_ASAP7_75t_R register___U12284 ( .A(register__n8089), .Y(register__n9721) );
  BUFx4f_ASAP7_75t_R register___U12285 ( .A(register__net106314), .Y(register__net101216) );
  BUFx2_ASAP7_75t_R register___U12286 ( .A(Reg_data[120]), .Y(register__net101217) );
  BUFx12f_ASAP7_75t_R register___U12287 ( .A(register__net89646), .Y(register__net89645) );
  BUFx6f_ASAP7_75t_R register___U12288 ( .A(register__net101216), .Y(register__net89646) );
  BUFx4f_ASAP7_75t_R register___U12289 ( .A(register__net134932), .Y(register__net101208) );
  BUFx2_ASAP7_75t_R register___U12290 ( .A(Reg_data[139]), .Y(register__net101209) );
  BUFx12f_ASAP7_75t_R register___U12291 ( .A(register__net88513), .Y(register__net88512) );
  BUFx6f_ASAP7_75t_R register___U12292 ( .A(register__net101208), .Y(register__net88513) );
  BUFx3_ASAP7_75t_R register___U12293 ( .A(register__n8093), .Y(register__n8092) );
  BUFx2_ASAP7_75t_R register___U12294 ( .A(Reg_data[348]), .Y(register__n8093) );
  BUFx4f_ASAP7_75t_R register___U12295 ( .A(register__net134033), .Y(register__net101198) );
  BUFx2_ASAP7_75t_R register___U12296 ( .A(Reg_data[189]), .Y(register__net101199) );
  BUFx6f_ASAP7_75t_R register___U12297 ( .A(register__net101198), .Y(register__net89566) );
  BUFx12f_ASAP7_75t_R register___U12298 ( .A(register__n8097), .Y(register__n8096) );
  BUFx12f_ASAP7_75t_R register___U12299 ( .A(register__n9522), .Y(register__n8097) );
  BUFx12f_ASAP7_75t_R register___U12300 ( .A(register__n8096), .Y(register__n9521) );
  BUFx6f_ASAP7_75t_R register___U12301 ( .A(register__n8094), .Y(register__n9522) );
  BUFx3_ASAP7_75t_R register___U12302 ( .A(register__n8099), .Y(register__n8098) );
  BUFx2_ASAP7_75t_R register___U12303 ( .A(Reg_data[375]), .Y(register__n8099) );
  BUFx3_ASAP7_75t_R register___U12304 ( .A(register__n8101), .Y(register__n8100) );
  BUFx2_ASAP7_75t_R register___U12305 ( .A(Reg_data[606]), .Y(register__n8101) );
  BUFx3_ASAP7_75t_R register___U12306 ( .A(register__n8103), .Y(register__n8102) );
  BUFx2_ASAP7_75t_R register___U12307 ( .A(Reg_data[365]), .Y(register__n8103) );
  BUFx2_ASAP7_75t_R register___U12308 ( .A(register__n9740), .Y(register__n8104) );
  BUFx2_ASAP7_75t_R register___U12309 ( .A(register__n9740), .Y(register__n8105) );
  BUFx4f_ASAP7_75t_R register___U12310 ( .A(register__n9740), .Y(register__n8106) );
  BUFx4f_ASAP7_75t_R register___U12311 ( .A(register__n6276), .Y(register__n8107) );
  BUFx2_ASAP7_75t_R register___U12312 ( .A(Reg_data[429]), .Y(register__n8108) );
  BUFx12f_ASAP7_75t_R register___U12313 ( .A(register__n9745), .Y(register__n8109) );
  BUFx12f_ASAP7_75t_R register___U12314 ( .A(register__n8109), .Y(register__n9744) );
  BUFx6f_ASAP7_75t_R register___U12315 ( .A(register__n8107), .Y(register__n9745) );
  BUFx4f_ASAP7_75t_R register___U12316 ( .A(register__n5831), .Y(register__n8110) );
  BUFx2_ASAP7_75t_R register___U12317 ( .A(Reg_data[941]), .Y(register__n8111) );
  BUFx12f_ASAP7_75t_R register___U12318 ( .A(register__n9755), .Y(register__n8112) );
  BUFx12f_ASAP7_75t_R register___U12319 ( .A(register__n8112), .Y(register__n9754) );
  BUFx6f_ASAP7_75t_R register___U12320 ( .A(register__n8110), .Y(register__n9755) );
  BUFx3_ASAP7_75t_R register___U12321 ( .A(register__n8114), .Y(register__n8113) );
  BUFx2_ASAP7_75t_R register___U12322 ( .A(Reg_data[141]), .Y(register__n8114) );
  BUFx4f_ASAP7_75t_R register___U12323 ( .A(register__n10146), .Y(register__n8115) );
  BUFx2_ASAP7_75t_R register___U12324 ( .A(register__n10146), .Y(register__n8116) );
  BUFx2_ASAP7_75t_R register___U12325 ( .A(register__n10146), .Y(register__n8117) );
  BUFx3_ASAP7_75t_R register___U12326 ( .A(register__n8119), .Y(register__n8118) );
  BUFx2_ASAP7_75t_R register___U12327 ( .A(Reg_data[173]), .Y(register__n8119) );
  BUFx12f_ASAP7_75t_R register___U12328 ( .A(register__n10149), .Y(register__n8120) );
  BUFx12f_ASAP7_75t_R register___U12329 ( .A(register__n8120), .Y(register__n10148) );
  BUFx2_ASAP7_75t_R register___U12330 ( .A(Reg_data[685]), .Y(register__n8122) );
  BUFx3_ASAP7_75t_R register___U12331 ( .A(register__net101127), .Y(register__net101126) );
  BUFx2_ASAP7_75t_R register___U12332 ( .A(Reg_data[157]), .Y(register__net101127) );
  BUFx3_ASAP7_75t_R register___U12333 ( .A(register__n8124), .Y(register__n8123) );
  BUFx2_ASAP7_75t_R register___U12334 ( .A(Reg_data[447]), .Y(register__n8124) );
  BUFx3_ASAP7_75t_R register___U12335 ( .A(register__n10503), .Y(register__n8125) );
  BUFx2_ASAP7_75t_R register___U12336 ( .A(register__n10503), .Y(register__n8126) );
  BUFx4f_ASAP7_75t_R register___U12337 ( .A(register__n10503), .Y(register__n8127) );
  BUFx3_ASAP7_75t_R register___U12338 ( .A(register__net101113), .Y(register__net101112) );
  BUFx2_ASAP7_75t_R register___U12339 ( .A(Reg_data[623]), .Y(register__net101113) );
  BUFx3_ASAP7_75t_R register___U12340 ( .A(register__n8129), .Y(register__n8128) );
  BUFx2_ASAP7_75t_R register___U12341 ( .A(Reg_data[218]), .Y(register__n8129) );
  BUFx3_ASAP7_75t_R register___U12342 ( .A(register__n8131), .Y(register__n8130) );
  BUFx2_ASAP7_75t_R register___U12343 ( .A(Reg_data[167]), .Y(register__n8131) );
  BUFx3_ASAP7_75t_R register___U12344 ( .A(register__n10179), .Y(register__n8132) );
  BUFx2_ASAP7_75t_R register___U12345 ( .A(register__n10179), .Y(register__n8133) );
  BUFx4f_ASAP7_75t_R register___U12346 ( .A(register__n10179), .Y(register__n8134) );
  BUFx3_ASAP7_75t_R register___U12347 ( .A(register__n8136), .Y(register__n8135) );
  BUFx2_ASAP7_75t_R register___U12348 ( .A(Reg_data[519]), .Y(register__n8136) );
  BUFx3_ASAP7_75t_R register___U12349 ( .A(register__n8138), .Y(register__n8137) );
  BUFx2_ASAP7_75t_R register___U12350 ( .A(Reg_data[604]), .Y(register__n8138) );
  BUFx3_ASAP7_75t_R register___U12351 ( .A(register__n8140), .Y(register__n8139) );
  BUFx2_ASAP7_75t_R register___U12352 ( .A(Reg_data[286]), .Y(register__n8140) );
  BUFx3_ASAP7_75t_R register___U12353 ( .A(register__n8142), .Y(register__n8141) );
  BUFx2_ASAP7_75t_R register___U12354 ( .A(Reg_data[830]), .Y(register__n8142) );
  BUFx3_ASAP7_75t_R register___U12355 ( .A(register__n8144), .Y(register__n8143) );
  BUFx2_ASAP7_75t_R register___U12356 ( .A(Reg_data[814]), .Y(register__n8144) );
  BUFx3_ASAP7_75t_R register___U12357 ( .A(register__n8146), .Y(register__n8145) );
  BUFx2_ASAP7_75t_R register___U12358 ( .A(Reg_data[926]), .Y(register__n8146) );
  BUFx2_ASAP7_75t_R register___U12359 ( .A(Reg_data[686]), .Y(register__n8148) );
  BUFx3_ASAP7_75t_R register___U12360 ( .A(register__n8150), .Y(register__n8149) );
  BUFx2_ASAP7_75t_R register___U12361 ( .A(Reg_data[785]), .Y(register__n8150) );
  BUFx4f_ASAP7_75t_R register___U12362 ( .A(register__net106297), .Y(register__net101055) );
  BUFx2_ASAP7_75t_R register___U12363 ( .A(Reg_data[874]), .Y(register__net101056) );
  BUFx12f_ASAP7_75t_R register___U12364 ( .A(register__net90458), .Y(register__net90457) );
  BUFx6f_ASAP7_75t_R register___U12365 ( .A(register__net101055), .Y(register__net90458) );
  BUFx3_ASAP7_75t_R register___U12366 ( .A(register__net101046), .Y(register__net101045) );
  BUFx2_ASAP7_75t_R register___U12367 ( .A(Reg_data[138]), .Y(register__net101046) );
  BUFx2_ASAP7_75t_R register___U12368 ( .A(register__net89289), .Y(register__net101048) );
  BUFx4f_ASAP7_75t_R register___U12369 ( .A(register__net89289), .Y(register__net101049) );
  BUFx3_ASAP7_75t_R register___U12370 ( .A(register__net101039), .Y(register__net101038) );
  BUFx2_ASAP7_75t_R register___U12371 ( .A(Reg_data[170]), .Y(register__net101039) );
  BUFx12f_ASAP7_75t_R register___U12372 ( .A(register__net89286), .Y(register__net89285) );
  BUFx3_ASAP7_75t_R register___U12373 ( .A(register__n8152), .Y(register__n8151) );
  BUFx2_ASAP7_75t_R register___U12374 ( .A(Reg_data[28]), .Y(register__n8152) );
  BUFx3_ASAP7_75t_R register___U12375 ( .A(register__n8154), .Y(register__n8153) );
  BUFx2_ASAP7_75t_R register___U12376 ( .A(Reg_data[140]), .Y(register__n8154) );
  BUFx4f_ASAP7_75t_R register___U12377 ( .A(register__n10225), .Y(register__n8155) );
  BUFx2_ASAP7_75t_R register___U12378 ( .A(register__n10225), .Y(register__n8156) );
  BUFx2_ASAP7_75t_R register___U12379 ( .A(register__n10225), .Y(register__n8157) );
  BUFx3_ASAP7_75t_R register___U12380 ( .A(register__n8159), .Y(register__n8158) );
  BUFx2_ASAP7_75t_R register___U12381 ( .A(Reg_data[819]), .Y(register__n8159) );
  BUFx2_ASAP7_75t_R register___U12382 ( .A(register__n9822), .Y(register__n8160) );
  BUFx2_ASAP7_75t_R register___U12383 ( .A(register__n9822), .Y(register__n8161) );
  BUFx4f_ASAP7_75t_R register___U12384 ( .A(register__n9822), .Y(register__n8162) );
  BUFx3_ASAP7_75t_R register___U12385 ( .A(register__n8164), .Y(register__n8163) );
  BUFx2_ASAP7_75t_R register___U12386 ( .A(Reg_data[147]), .Y(register__n8164) );
  BUFx3_ASAP7_75t_R register___U12387 ( .A(register__net101001), .Y(register__net101000) );
  BUFx2_ASAP7_75t_R register___U12388 ( .A(Reg_data[394]), .Y(register__net101001) );
  BUFx2_ASAP7_75t_R register___U12389 ( .A(register__net90397), .Y(register__net101003) );
  BUFx4f_ASAP7_75t_R register___U12390 ( .A(register__net90397), .Y(register__net101004) );
  BUFx3_ASAP7_75t_R register___U12391 ( .A(register__net100991), .Y(register__net100990) );
  BUFx2_ASAP7_75t_R register___U12392 ( .A(Reg_data[42]), .Y(register__net100991) );
  BUFx4f_ASAP7_75t_R register___U12393 ( .A(register__net89213), .Y(register__net100992) );
  BUFx2_ASAP7_75t_R register___U12394 ( .A(register__net89213), .Y(register__net100994) );
  BUFx2_ASAP7_75t_R register___U12395 ( .A(Reg_data[955]), .Y(register__n8166) );
  BUFx3_ASAP7_75t_R register___U12396 ( .A(register__n8168), .Y(register__n8167) );
  BUFx2_ASAP7_75t_R register___U12397 ( .A(Reg_data[155]), .Y(register__n8168) );
  BUFx3_ASAP7_75t_R register___U12398 ( .A(register__n10265), .Y(register__n8169) );
  BUFx2_ASAP7_75t_R register___U12399 ( .A(register__n10265), .Y(register__n8170) );
  BUFx4f_ASAP7_75t_R register___U12400 ( .A(register__n10265), .Y(register__n8171) );
  BUFx2_ASAP7_75t_R register___U12401 ( .A(Reg_data[55]), .Y(register__n8173) );
  BUFx3_ASAP7_75t_R register___U12402 ( .A(register__n8175), .Y(register__n8174) );
  BUFx2_ASAP7_75t_R register___U12403 ( .A(Reg_data[361]), .Y(register__n8175) );
  BUFx3_ASAP7_75t_R register___U12404 ( .A(register__n8177), .Y(register__n8176) );
  BUFx2_ASAP7_75t_R register___U12405 ( .A(Reg_data[41]), .Y(register__n8177) );
  BUFx12f_ASAP7_75t_R register___U12406 ( .A(register__n10274), .Y(register__n8178) );
  BUFx12f_ASAP7_75t_R register___U12407 ( .A(register__n8178), .Y(register__n10273) );
  BUFx4f_ASAP7_75t_R register___U12408 ( .A(register__n6279), .Y(register__n8179) );
  BUFx2_ASAP7_75t_R register___U12409 ( .A(Reg_data[826]), .Y(register__n8180) );
  BUFx12f_ASAP7_75t_R register___U12410 ( .A(register__n9854), .Y(register__n8181) );
  BUFx12f_ASAP7_75t_R register___U12411 ( .A(register__n8181), .Y(register__n9853) );
  BUFx6f_ASAP7_75t_R register___U12412 ( .A(register__n8179), .Y(register__n9854) );
  BUFx4f_ASAP7_75t_R register___U12413 ( .A(register__n5178), .Y(register__n8182) );
  BUFx2_ASAP7_75t_R register___U12414 ( .A(Reg_data[954]), .Y(register__n8183) );
  BUFx12f_ASAP7_75t_R register___U12415 ( .A(register__n9856), .Y(register__n9855) );
  BUFx6f_ASAP7_75t_R register___U12416 ( .A(register__n8182), .Y(register__n9856) );
  BUFx3_ASAP7_75t_R register___U12417 ( .A(register__n8185), .Y(register__n8184) );
  BUFx2_ASAP7_75t_R register___U12418 ( .A(Reg_data[186]), .Y(register__n8185) );
  BUFx12f_ASAP7_75t_R register___U12419 ( .A(register__n10282), .Y(register__n8186) );
  BUFx12f_ASAP7_75t_R register___U12420 ( .A(register__n8186), .Y(register__n10281) );
  BUFx3_ASAP7_75t_R register___U12421 ( .A(register__n8188), .Y(register__n8187) );
  BUFx2_ASAP7_75t_R register___U12422 ( .A(Reg_data[767]), .Y(register__n8188) );
  BUFx12f_ASAP7_75t_R register___U12423 ( .A(register__n5659), .Y(register__n8779) );
  BUFx4f_ASAP7_75t_R register___U12424 ( .A(register__n6535), .Y(register__n8189) );
  BUFx2_ASAP7_75t_R register___U12425 ( .A(Reg_data[959]), .Y(register__n8190) );
  BUFx12f_ASAP7_75t_R register___U12426 ( .A(register__n9862), .Y(register__n9861) );
  BUFx6f_ASAP7_75t_R register___U12427 ( .A(register__n8189), .Y(register__n9862) );
  BUFx3_ASAP7_75t_R register___U12428 ( .A(register__n8192), .Y(register__n8191) );
  BUFx2_ASAP7_75t_R register___U12429 ( .A(Reg_data[364]), .Y(register__n8192) );
  BUFx3_ASAP7_75t_R register___U12430 ( .A(register__n9875), .Y(register__n8193) );
  BUFx6f_ASAP7_75t_R register___U12431 ( .A(register__n9875), .Y(register__n8194) );
  BUFx3_ASAP7_75t_R register___U12432 ( .A(register__n8196), .Y(register__n8195) );
  BUFx2_ASAP7_75t_R register___U12433 ( .A(Reg_data[433]), .Y(register__n8196) );
  BUFx12f_ASAP7_75t_R register___U12434 ( .A(register__n9888), .Y(register__n8197) );
  BUFx12f_ASAP7_75t_R register___U12435 ( .A(register__n8197), .Y(register__n9887) );
  BUFx4f_ASAP7_75t_R register___U12436 ( .A(register__net118011), .Y(register__net100902) );
  BUFx2_ASAP7_75t_R register___U12437 ( .A(Reg_data[952]), .Y(register__net100903) );
  BUFx6f_ASAP7_75t_R register___U12438 ( .A(register__net100902), .Y(register__net90249) );
  BUFx3_ASAP7_75t_R register___U12439 ( .A(register__net100893), .Y(register__net100892) );
  BUFx2_ASAP7_75t_R register___U12440 ( .A(Reg_data[152]), .Y(register__net100893) );
  BUFx4f_ASAP7_75t_R register___U12441 ( .A(register__net89053), .Y(register__net100894) );
  BUFx2_ASAP7_75t_R register___U12442 ( .A(register__net89053), .Y(register__net100896) );
  BUFx3_ASAP7_75t_R register___U12443 ( .A(register__net100886), .Y(register__net100885) );
  BUFx2_ASAP7_75t_R register___U12444 ( .A(Reg_data[184]), .Y(register__net100886) );
  BUFx12f_ASAP7_75t_R register___U12445 ( .A(register__net89050), .Y(register__net89049) );
  BUFx3_ASAP7_75t_R register___U12446 ( .A(register__n8199), .Y(register__n8198) );
  BUFx2_ASAP7_75t_R register___U12447 ( .A(Reg_data[219]), .Y(register__n8199) );
  BUFx3_ASAP7_75t_R register___U12448 ( .A(register__n10513), .Y(register__n8200) );
  BUFx2_ASAP7_75t_R register___U12449 ( .A(register__n10513), .Y(register__n8201) );
  BUFx3_ASAP7_75t_R register___U12450 ( .A(register__n8204), .Y(register__n8203) );
  BUFx2_ASAP7_75t_R register___U12451 ( .A(Reg_data[924]), .Y(register__n8204) );
  BUFx3_ASAP7_75t_R register___U12452 ( .A(register__n9899), .Y(register__n8205) );
  BUFx2_ASAP7_75t_R register___U12453 ( .A(register__n9899), .Y(register__n8206) );
  BUFx4f_ASAP7_75t_R register___U12454 ( .A(register__n9899), .Y(register__n8207) );
  BUFx3_ASAP7_75t_R register___U12455 ( .A(register__n8209), .Y(register__n8208) );
  BUFx2_ASAP7_75t_R register___U12456 ( .A(Reg_data[700]), .Y(register__n8209) );
  BUFx4f_ASAP7_75t_R register___U12457 ( .A(register__n7712), .Y(register__n8210) );
  BUFx12f_ASAP7_75t_R register___U12458 ( .A(register__n8213), .Y(register__n8212) );
  BUFx12f_ASAP7_75t_R register___U12459 ( .A(register__n10420), .Y(register__n8213) );
  BUFx12f_ASAP7_75t_R register___U12460 ( .A(register__n8212), .Y(register__n10419) );
  BUFx6f_ASAP7_75t_R register___U12461 ( .A(register__n8210), .Y(register__n10420) );
  BUFx3_ASAP7_75t_R register___U12462 ( .A(register__n8215), .Y(register__n8214) );
  BUFx2_ASAP7_75t_R register___U12463 ( .A(Reg_data[732]), .Y(register__n8215) );
  BUFx4f_ASAP7_75t_R register___U12464 ( .A(register__n11436), .Y(register__n8216) );
  INVx2_ASAP7_75t_R register___U12465 ( .A(register__n8718), .Y(register__n11436) );
  BUFx6f_ASAP7_75t_R register___U12466 ( .A(register__n8719), .Y(register__n8718) );
  INVx2_ASAP7_75t_R register___U12467 ( .A(register__net97197), .Y(register__net100833) );
  BUFx6f_ASAP7_75t_R register___U12468 ( .A(register__net97198), .Y(register__net97197) );
  BUFx12f_ASAP7_75t_R register___U12469 ( .A(register__net62712), .Y(register__net100796) );
  BUFx12f_ASAP7_75t_R register___U12470 ( .A(register__net100799), .Y(register__net100797) );
  BUFx12f_ASAP7_75t_R register___U12471 ( .A(register__net143790), .Y(register__net62706) );
  INVx1_ASAP7_75t_R register___U12472 ( .A(register__n5284), .Y(register__n8217) );
  INVx1_ASAP7_75t_R register___U12473 ( .A(register__n5591), .Y(register__n8218) );
  INVx1_ASAP7_75t_R register___U12474 ( .A(register__n5593), .Y(register__n8219) );
  INVx1_ASAP7_75t_R register___U12475 ( .A(register__n5595), .Y(register__n8220) );
  INVx1_ASAP7_75t_R register___U12476 ( .A(register__n4801), .Y(register__n8222) );
  INVx1_ASAP7_75t_R register___U12477 ( .A(register__n4803), .Y(register__n8223) );
  INVx1_ASAP7_75t_R register___U12478 ( .A(register__n4805), .Y(register__n8224) );
  INVx1_ASAP7_75t_R register___U12479 ( .A(register__n10905), .Y(register__n8228) );
  AO22x1_ASAP7_75t_R register___U12480 ( .A1(register__n8515), .A2(register__C6423_net61318), .B1(register__n6661), 
        .B2(register__n1446), .Y(register__n11628) );
  INVx1_ASAP7_75t_R register___U12481 ( .A(register__n4738), .Y(register__n8229) );
  INVx1_ASAP7_75t_R register___U12482 ( .A(register__n3207), .Y(register__n8230) );
  INVx1_ASAP7_75t_R register___U12483 ( .A(register__n4173), .Y(register__n8231) );
  INVx1_ASAP7_75t_R register___U12484 ( .A(register__n4175), .Y(register__n8232) );
  INVx1_ASAP7_75t_R register___U12485 ( .A(register__n11012), .Y(register__n8234) );
  INVx1_ASAP7_75t_R register___U12486 ( .A(register__n5253), .Y(register__n8235) );
  INVx1_ASAP7_75t_R register___U12487 ( .A(register__n10731), .Y(register__n8236) );
  BUFx6f_ASAP7_75t_R register___U12488 ( .A(register__net100610), .Y(register__net63374) );
  BUFx6f_ASAP7_75t_R register___U12489 ( .A(register__net100610), .Y(register__net63376) );
  BUFx6f_ASAP7_75t_R register___U12490 ( .A(register__net100610), .Y(register__net63368) );
  BUFx6f_ASAP7_75t_R register___U12491 ( .A(register__net100610), .Y(register__net63370) );
  OA22x2_ASAP7_75t_R register___U12492 ( .A1(register__n12225), .A2(register__n1988), .B1(register__n10120), .B2(register__n3170), 
        .Y(register__n13346) );
  OA22x2_ASAP7_75t_R register___U12493 ( .A1(register__n11949), .A2(register__n1988), .B1(register__n10458), .B2(register__n11734), .Y(register__n13356) );
  OA22x2_ASAP7_75t_R register___U12494 ( .A1(register__n12142), .A2(register__n1988), .B1(register__n10102), .B2(register__n3267), 
        .Y(register__n13349) );
  OA22x2_ASAP7_75t_R register___U12495 ( .A1(register__n3700), .A2(register__n1001), .B1(register__n10068), .B2(register__n970), 
        .Y(register__n13206) );
  INVx1_ASAP7_75t_R register___U12496 ( .A(register__n3895), .Y(register__n8237) );
  OA22x2_ASAP7_75t_R register___U12497 ( .A1(register__n12367), .A2(register__n991), .B1(register__n10076), .B2(register__n969), 
        .Y(register__n13186) );
  OA22x2_ASAP7_75t_R register___U12498 ( .A1(register__net64754), .A2(register__n987), .B1(register__net89689), .B2(
        n972), .Y(register__n13202) );
  OA22x2_ASAP7_75t_R register___U12499 ( .A1(register__net64922), .A2(register__n990), .B1(register__n10091), .B2(register__n974), 
        .Y(register__n13204) );
  INVx1_ASAP7_75t_R register___U12500 ( .A(register__n6246), .Y(register__n8239) );
  OA22x2_ASAP7_75t_R register___U12501 ( .A1(register__net63236), .A2(register__n1989), .B1(register__net89421), .B2(
        n3392), .Y(register__n13340) );
  OA22x2_ASAP7_75t_R register___U12502 ( .A1(register__net63242), .A2(register__n993), .B1(register__net89413), .B2(
        n971), .Y(register__n13184) );
  INVx1_ASAP7_75t_R register___U12503 ( .A(register__n5977), .Y(register__n8241) );
  INVx1_ASAP7_75t_R register___U12504 ( .A(register__n5979), .Y(register__n8242) );
  OA22x2_ASAP7_75t_R register___U12505 ( .A1(register__net62654), .A2(register__n1000), .B1(register__n9371), .B2(register__n971), 
        .Y(register__n13177) );
  INVx1_ASAP7_75t_R register___U12506 ( .A(register__n6258), .Y(register__n8243) );
  OA22x2_ASAP7_75t_R register___U12507 ( .A1(register__n12453), .A2(register__n2851), .B1(register__n10199), .B2(register__n11747), .Y(register__n13263) );
  OA22x2_ASAP7_75t_R register___U12508 ( .A1(register__n12420), .A2(register__n1988), .B1(register__n9369), .B2(register__n5183), 
        .Y(register__n13337) );
  BUFx6f_ASAP7_75t_R register___U12509 ( .A(register__net100539), .Y(register__net64466) );
  BUFx12f_ASAP7_75t_R register___U12510 ( .A(register__net100542), .Y(register__net64464) );
  BUFx16f_ASAP7_75t_R register___U12511 ( .A(register__net137769), .Y(register__net64474) );
  BUFx6f_ASAP7_75t_R register___U12512 ( .A(register__n4835), .Y(register__n12328) );
  BUFx6f_ASAP7_75t_R register___U12513 ( .A(register__n12329), .Y(register__n12324) );
  BUFx2_ASAP7_75t_R register___U12514 ( .A(register__n12334), .Y(register__n12327) );
  BUFx6f_ASAP7_75t_R register___U12515 ( .A(register__n3533), .Y(register__n12270) );
  BUFx6f_ASAP7_75t_R register___U12516 ( .A(register__n4576), .Y(register__n12275) );
  BUFx6f_ASAP7_75t_R register___U12517 ( .A(register__n12098), .Y(register__n12099) );
  BUFx6f_ASAP7_75t_R register___U12518 ( .A(register__n5041), .Y(register__n12187) );
  BUFx6f_ASAP7_75t_R register___U12519 ( .A(register__n3677), .Y(register__n12186) );
  INVx1_ASAP7_75t_R register___U12520 ( .A(register__n5613), .Y(register__n8251) );
  INVx1_ASAP7_75t_R register___U12521 ( .A(register__n4688), .Y(register__n8252) );
  INVx1_ASAP7_75t_R register___U12522 ( .A(register__n4690), .Y(register__n8253) );
  INVx1_ASAP7_75t_R register___U12523 ( .A(register__n4692), .Y(register__n8254) );
  INVx1_ASAP7_75t_R register___U12524 ( .A(register__n5555), .Y(register__n8256) );
  INVx1_ASAP7_75t_R register___U12525 ( .A(register__n4547), .Y(register__n8258) );
  INVx1_ASAP7_75t_R register___U12526 ( .A(register__n4549), .Y(register__n8259) );
  INVx1_ASAP7_75t_R register___U12527 ( .A(register__n4905), .Y(register__n8262) );
  INVx1_ASAP7_75t_R register___U12528 ( .A(register__n11120), .Y(register__n8264) );
  INVx1_ASAP7_75t_R register___U12529 ( .A(register__n4441), .Y(register__n8266) );
  INVx1_ASAP7_75t_R register___U12530 ( .A(register__n4627), .Y(register__n8269) );
  INVx1_ASAP7_75t_R register___U12531 ( .A(register__n4629), .Y(register__n8270) );
  INVx1_ASAP7_75t_R register___U12532 ( .A(register__n4743), .Y(register__n8274) );
  INVx1_ASAP7_75t_R register___U12533 ( .A(register__n3166), .Y(register__n8275) );
  INVx1_ASAP7_75t_R register___U12534 ( .A(register__n5616), .Y(register__n8276) );
  INVx4_ASAP7_75t_R register___U12535 ( .A(register__net62710), .Y(register__net62674) );
  OA22x2_ASAP7_75t_R register___U12536 ( .A1(register__n12345), .A2(register__n1988), .B1(register__n10074), .B2(register__n3391), 
        .Y(register__n13342) );
  OA22x2_ASAP7_75t_R register___U12537 ( .A1(register__n12279), .A2(register__n1989), .B1(register__n10158), .B2(register__n3390), 
        .Y(register__n13344) );
  OA22x2_ASAP7_75t_R register___U12538 ( .A1(register__n12405), .A2(register__n997), .B1(register__n10165), .B2(register__n970), 
        .Y(register__n13182) );
  INVx1_ASAP7_75t_R register___U12539 ( .A(register__n6793), .Y(register__n8280) );
  OA22x2_ASAP7_75t_R register___U12540 ( .A1(register__n3319), .A2(register__n995), .B1(register__n10153), .B2(register__n969), 
        .Y(register__n13180) );
  INVx1_ASAP7_75t_R register___U12541 ( .A(register__n4409), .Y(register__n8281) );
  INVx2_ASAP7_75t_R register___U12542 ( .A(register__n12439), .Y(register__n12423) );
  OA22x2_ASAP7_75t_R register___U12543 ( .A1(register__n12421), .A2(register__n701), .B1(register__n10393), .B2(register__n672), 
        .Y(register__n13309) );
  OR3x1_ASAP7_75t_R register___U12544 ( .A(register__n5323), .B(register__n8286), .C(register__n8285), .Y(register__n11475) );
  OA22x2_ASAP7_75t_R register___U12545 ( .A1(register__net131654), .A2(register__n6768), .B1(register__net130175), .B2(
        n10867), .Y(register__n11478) );
  OA22x2_ASAP7_75t_R register___U12546 ( .A1(register__n710), .A2(register__n7870), .B1(register__n1113), .B2(register__n7091), 
        .Y(register__n11477) );
  INVx1_ASAP7_75t_R register___U12547 ( .A(register__n5321), .Y(register__n8286) );
  OA222x2_ASAP7_75t_R register___U12548 ( .A1(register__n1987), .A2(register__n10870), .B1(register__n1995), .B2(register__n7579), 
        .C1(register__n1800), .C2(register__n6205), .Y(register__n11476) );
  OR3x1_ASAP7_75t_R register___U12549 ( .A(register__n5144), .B(register__n8288), .C(register__n8287), .Y(register__n10700) );
  OA22x2_ASAP7_75t_R register___U12550 ( .A1(register__n419), .A2(register__net113227), .B1(register__n800), .B2(
        net103295), .Y(register__n10703) );
  INVx1_ASAP7_75t_R register___U12551 ( .A(register__n5140), .Y(register__n8287) );
  OA22x2_ASAP7_75t_R register___U12552 ( .A1(register__net107674), .A2(register__C6423_net60749), .B1(register__n1691), 
        .B2(register__C6422_net59832), .Y(register__n10702) );
  INVx1_ASAP7_75t_R register___U12553 ( .A(register__n5142), .Y(register__n8288) );
  OA222x2_ASAP7_75t_R register___U12554 ( .A1(register__n2002), .A2(register__net115136), .B1(register__n817), .B2(
        net105530), .C1(register__net112580), .C2(register__C6422_net59835), .Y(register__n10701) );
  OR3x1_ASAP7_75t_R register___U12555 ( .A(register__n773), .B(register__n8290), .C(register__n2228), .Y(register__n11344) );
  OA22x2_ASAP7_75t_R register___U12556 ( .A1(register__net131654), .A2(register__n7689), .B1(register__net130175), .B2(
        n8589), .Y(register__n11347) );
  OA22x2_ASAP7_75t_R register___U12557 ( .A1(register__n711), .A2(register__n7100), .B1(register__n353), .B2(register__n7582), 
        .Y(register__n11346) );
  INVx1_ASAP7_75t_R register___U12558 ( .A(register__n6008), .Y(register__n8290) );
  OA222x2_ASAP7_75t_R register___U12559 ( .A1(register__n1987), .A2(register__n6476), .B1(register__n1995), .B2(register__n5726), 
        .C1(register__n1800), .C2(register__n6213), .Y(register__n11345) );
  OR3x1_ASAP7_75t_R register___U12560 ( .A(register__n5466), .B(register__n8293), .C(register__n8292), .Y(register__n10886) );
  OA22x2_ASAP7_75t_R register___U12561 ( .A1(register__n420), .A2(register__n7101), .B1(register__n802), .B2(register__n8591), 
        .Y(register__n10889) );
  INVx1_ASAP7_75t_R register___U12562 ( .A(register__n5462), .Y(register__n8292) );
  OA22x2_ASAP7_75t_R register___U12563 ( .A1(register__net107674), .A2(register__n11501), .B1(register__n1691), .B2(
        n7583), .Y(register__n10888) );
  INVx1_ASAP7_75t_R register___U12564 ( .A(register__n5464), .Y(register__n8293) );
  OA222x2_ASAP7_75t_R register___U12565 ( .A1(register__n2081), .A2(register__n6223), .B1(register__n817), .B2(register__n11503), 
        .C1(register__net112578), .C2(register__n6471), .Y(register__n10887) );
  INVx1_ASAP7_75t_R register___U12566 ( .A(register__n10887), .Y(register__n8294) );
  OR3x1_ASAP7_75t_R register___U12567 ( .A(register__n5493), .B(register__n8297), .C(register__n8296), .Y(register__n11081) );
  OA22x2_ASAP7_75t_R register___U12568 ( .A1(register__n420), .A2(register__C6422_net60323), .B1(register__n801), .B2(
        C6422_net60324), .Y(register__n11084) );
  INVx1_ASAP7_75t_R register___U12569 ( .A(register__n5489), .Y(register__n8296) );
  OA22x2_ASAP7_75t_R register___U12570 ( .A1(register__net107674), .A2(register__net105488), .B1(register__n1691), .B2(
        net108748), .Y(register__n11083) );
  INVx1_ASAP7_75t_R register___U12571 ( .A(register__n5491), .Y(register__n8297) );
  OA222x2_ASAP7_75t_R register___U12572 ( .A1(register__n2002), .A2(register__C6423_net61245), .B1(register__n817), 
        .B2(register__C6422_net60328), .C1(register__net112580), .C2(register__C6422_net60329), .Y(register__n11082)
         );
  INVx1_ASAP7_75t_R register___U12573 ( .A(register__n11082), .Y(register__n8298) );
  OR3x1_ASAP7_75t_R register___U12574 ( .A(register__n5805), .B(register__n8300), .C(register__n8299), .Y(register__n11520) );
  OA22x2_ASAP7_75t_R register___U12575 ( .A1(register__n2013), .A2(register__n6767), .B1(register__net130175), .B2(
        n10914), .Y(register__n11523) );
  INVx1_ASAP7_75t_R register___U12576 ( .A(register__n11523), .Y(register__n8299) );
  OR3x1_ASAP7_75t_R register___U12577 ( .A(register__n5129), .B(register__n8304), .C(register__n8303), .Y(register__n10525) );
  OA22x2_ASAP7_75t_R register___U12578 ( .A1(register__n419), .A2(register__n7094), .B1(register__n800), .B2(register__n6228), 
        .Y(register__n10528) );
  OA22x2_ASAP7_75t_R register___U12579 ( .A1(register__net107674), .A2(register__n7869), .B1(register__n1691), .B2(
        n6765), .Y(register__n10527) );
  INVx1_ASAP7_75t_R register___U12580 ( .A(register__n5126), .Y(register__n8304) );
  OR3x1_ASAP7_75t_R register___U12581 ( .A(register__n4828), .B(register__n8307), .C(register__n8306), .Y(register__n10614) );
  OA22x2_ASAP7_75t_R register___U12582 ( .A1(register__n420), .A2(register__n10618), .B1(register__n802), .B2(register__n6985), 
        .Y(register__n10617) );
  INVx1_ASAP7_75t_R register___U12583 ( .A(register__n4824), .Y(register__n8306) );
  OA22x2_ASAP7_75t_R register___U12584 ( .A1(register__net107674), .A2(register__n7586), .B1(register__n1691), .B2(
        n7243), .Y(register__n10616) );
  INVx1_ASAP7_75t_R register___U12585 ( .A(register__n4826), .Y(register__n8307) );
  INVx1_ASAP7_75t_R register___U12586 ( .A(register__n10615), .Y(register__n8308) );
  OR3x1_ASAP7_75t_R register___U12587 ( .A(register__n4946), .B(register__n8310), .C(register__n8309), .Y(register__n10636) );
  OA22x2_ASAP7_75t_R register___U12588 ( .A1(register__n420), .A2(register__n8837), .B1(register__n800), .B2(register__n11305), 
        .Y(register__n10638) );
  INVx1_ASAP7_75t_R register___U12589 ( .A(register__n4944), .Y(register__n8309) );
  OA22x2_ASAP7_75t_R register___U12590 ( .A1(register__net107674), .A2(register__n9148), .B1(register__n1691), .B2(
        n7245), .Y(register__n10637) );
  OR3x1_ASAP7_75t_R register___U12591 ( .A(register__n5161), .B(register__n8313), .C(register__n8311), .Y(register__n10802) );
  OA22x2_ASAP7_75t_R register___U12592 ( .A1(register__n419), .A2(register__net108770), .B1(register__n800), .B2(
        net113150), .Y(register__n10805) );
  INVx1_ASAP7_75t_R register___U12593 ( .A(register__n5158), .Y(register__n8311) );
  OA22x2_ASAP7_75t_R register___U12594 ( .A1(register__n66), .A2(register__C6422_net59961), .B1(register__n1691), .B2(
        C6423_net60880), .Y(register__n10804) );
  INVx1_ASAP7_75t_R register___U12595 ( .A(register__n5162), .Y(register__n8313) );
  OR3x1_ASAP7_75t_R register___U12596 ( .A(register__n364), .B(register__n8316), .C(register__n8315), .Y(register__n10929) );
  OA22x2_ASAP7_75t_R register___U12597 ( .A1(register__n420), .A2(register__n6771), .B1(register__n800), .B2(register__n6480), 
        .Y(register__n10932) );
  INVx1_ASAP7_75t_R register___U12598 ( .A(register__n4935), .Y(register__n8315) );
  OA22x2_ASAP7_75t_R register___U12599 ( .A1(register__net107674), .A2(register__n6229), .B1(register__n1691), .B2(
        n7095), .Y(register__n10931) );
  INVx1_ASAP7_75t_R register___U12600 ( .A(register__n4937), .Y(register__n8316) );
  OA222x2_ASAP7_75t_R register___U12601 ( .A1(register__n1978), .A2(register__n11547), .B1(register__n1117), .B2(register__n7581), 
        .C1(register__net112580), .C2(register__n7866), .Y(register__n10930) );
  OR3x1_ASAP7_75t_R register___U12602 ( .A(register__n5470), .B(register__n8318), .C(register__n8317), .Y(register__n10735) );
  OA22x2_ASAP7_75t_R register___U12603 ( .A1(register__n420), .A2(register__n7102), .B1(register__n800), .B2(register__n8590), 
        .Y(register__n10738) );
  INVx1_ASAP7_75t_R register___U12604 ( .A(register__n5467), .Y(register__n8317) );
  OA22x2_ASAP7_75t_R register___U12605 ( .A1(register__n66), .A2(register__n7694), .B1(register__n1691), .B2(register__n11372), 
        .Y(register__n10737) );
  OA222x2_ASAP7_75t_R register___U12606 ( .A1(register__n2002), .A2(register__n6224), .B1(register__n817), .B2(register__n5727), 
        .C1(register__net112580), .C2(register__n7578), .Y(register__n10736) );
  INVx1_ASAP7_75t_R register___U12607 ( .A(register__n5469), .Y(register__n8319) );
  OR3x1_ASAP7_75t_R register___U12608 ( .A(register__n5340), .B(register__n8321), .C(register__n8320), .Y(register__n11701) );
  OA22x2_ASAP7_75t_R register___U12609 ( .A1(register__net131654), .A2(register__n11705), .B1(register__net130175), 
        .B2(register__n11706), .Y(register__n11704) );
  INVx1_ASAP7_75t_R register___U12610 ( .A(register__n5338), .Y(register__n8320) );
  OA22x2_ASAP7_75t_R register___U12611 ( .A1(register__n714), .A2(register__n7104), .B1(register__net149933), .B2(
        n11129), .Y(register__n11703) );
  INVx1_ASAP7_75t_R register___U12612 ( .A(register__n5339), .Y(register__n8321) );
  OR3x1_ASAP7_75t_R register___U12613 ( .A(register__n5169), .B(register__n8324), .C(register__n8323), .Y(register__n11013) );
  OA22x2_ASAP7_75t_R register___U12614 ( .A1(register__n420), .A2(register__n6490), .B1(register__n800), .B2(register__n9159), 
        .Y(register__n11016) );
  INVx1_ASAP7_75t_R register___U12615 ( .A(register__n5163), .Y(register__n8323) );
  OA22x2_ASAP7_75t_R register___U12616 ( .A1(register__net107674), .A2(register__n8363), .B1(register__n1691), .B2(
        n7108), .Y(register__n11015) );
  INVx1_ASAP7_75t_R register___U12617 ( .A(register__n5165), .Y(register__n8324) );
  OA222x2_ASAP7_75t_R register___U12618 ( .A1(register__n2002), .A2(register__n6226), .B1(register__n817), .B2(register__n5955), 
        .C1(register__net112580), .C2(register__n7577), .Y(register__n11014) );
  OA22x2_ASAP7_75t_R register___U12619 ( .A1(register__n1964), .A2(register__n8361), .B1(register__net130175), .B2(
        n7346), .Y(register__n11642) );
  INVx1_ASAP7_75t_R register___U12620 ( .A(register__n6028), .Y(register__n8326) );
  OA222x2_ASAP7_75t_R register___U12621 ( .A1(register__n1987), .A2(register__n11043), .B1(register__n1995), .B2(
        net108812), .C1(register__n1800), .C2(register__net103310), .Y(register__n11641) );
  INVx3_ASAP7_75t_R register___U12622 ( .A(register__n7717), .Y(register__n11645) );
  INVx3_ASAP7_75t_R register___U12623 ( .A(register__n7720), .Y(register__n11042) );
  BUFx12f_ASAP7_75t_R register___U12624 ( .A(register__n3606), .Y(register__n8334) );
  BUFx12f_ASAP7_75t_R register___U12625 ( .A(register__n11743), .Y(register__n8336) );
  OA22x2_ASAP7_75t_R register___U12626 ( .A1(register__net131654), .A2(register__n7103), .B1(register__net130175), .B2(
        n7868), .Y(register__n11411) );
  INVx1_ASAP7_75t_R register___U12627 ( .A(register__n5820), .Y(register__n8339) );
  OA22x2_ASAP7_75t_R register___U12628 ( .A1(register__n710), .A2(register__n6764), .B1(register__n1113), .B2(register__n7584), 
        .Y(register__n11410) );
  INVx1_ASAP7_75t_R register___U12629 ( .A(register__n5822), .Y(register__n8340) );
  OA222x2_ASAP7_75t_R register___U12630 ( .A1(register__n1987), .A2(register__n6225), .B1(register__n1995), .B2(register__n6472), 
        .C1(register__n1800), .C2(register__n10789), .Y(register__n11409) );
  BUFx6f_ASAP7_75t_R register___U12631 ( .A(register__n8342), .Y(register__n8341) );
  BUFx4f_ASAP7_75t_R register___U12632 ( .A(register__n5195), .Y(register__n8342) );
  BUFx6f_ASAP7_75t_R register___U12633 ( .A(register__n8344), .Y(register__n8343) );
  BUFx4f_ASAP7_75t_R register___U12634 ( .A(register__n7404), .Y(register__n8344) );
  BUFx6f_ASAP7_75t_R register___U12635 ( .A(register__n8346), .Y(register__n8345) );
  BUFx4f_ASAP7_75t_R register___U12636 ( .A(register__n6070), .Y(register__n8346) );
  BUFx6f_ASAP7_75t_R register___U12637 ( .A(register__n8350), .Y(register__n8349) );
  BUFx4f_ASAP7_75t_R register___U12638 ( .A(register__n6589), .Y(register__n8350) );
  BUFx4f_ASAP7_75t_R register___U12639 ( .A(register__n7541), .Y(register__n8352) );
  BUFx6f_ASAP7_75t_R register___U12640 ( .A(register__n8355), .Y(register__n8354) );
  BUFx4f_ASAP7_75t_R register___U12641 ( .A(register__n6390), .Y(register__n8355) );
  BUFx6f_ASAP7_75t_R register___U12642 ( .A(register__n8357), .Y(register__n8356) );
  BUFx4f_ASAP7_75t_R register___U12643 ( .A(register__n6622), .Y(register__n8357) );
  INVx2_ASAP7_75t_R register___U12644 ( .A(register__n11736), .Y(register__n11854) );
  BUFx2_ASAP7_75t_R register___U12645 ( .A(register__n11327), .Y(register__n8359) );
  BUFx2_ASAP7_75t_R register___U12646 ( .A(register__n10661), .Y(register__n8360) );
  BUFx2_ASAP7_75t_R register___U12647 ( .A(register__C6423_net61111), .Y(register__net99209) );
  BUFx2_ASAP7_75t_R register___U12648 ( .A(register__n11643), .Y(register__n8361) );
  BUFx2_ASAP7_75t_R register___U12649 ( .A(register__n11305), .Y(register__n8362) );
  BUFx2_ASAP7_75t_R register___U12650 ( .A(register__n11018), .Y(register__n8363) );
  BUFx2_ASAP7_75t_R register___U12651 ( .A(register__n12931), .Y(register__n8365) );
  BUFx2_ASAP7_75t_R register___U12652 ( .A(register__n8367), .Y(register__n8366) );
  BUFx2_ASAP7_75t_R register___U12653 ( .A(register__n13061), .Y(register__n8367) );
  INVx3_ASAP7_75t_R register___U12654 ( .A(register__n12445), .Y(register__n12429) );
  BUFx6f_ASAP7_75t_R register___U12655 ( .A(register__net99038), .Y(register__net99037) );
  BUFx4f_ASAP7_75t_R register___U12656 ( .A(register__C6423_net60878), .Y(register__net99038) );
  BUFx6f_ASAP7_75t_R register___U12657 ( .A(register__net99034), .Y(register__net99033) );
  BUFx4f_ASAP7_75t_R register___U12658 ( .A(register__C6423_net61090), .Y(register__net99034) );
  BUFx12f_ASAP7_75t_R register___U12659 ( .A(register__n9707), .Y(register__n8368) );
  BUFx3_ASAP7_75t_R register___U12660 ( .A(register__n8938), .Y(register__n8369) );
  BUFx3_ASAP7_75t_R register___U12661 ( .A(register__n8987), .Y(register__n8371) );
  BUFx4f_ASAP7_75t_R register___U12662 ( .A(register__net90677), .Y(register__net95244) );
  BUFx3_ASAP7_75t_R register___U12663 ( .A(register__net95809), .Y(register__net98937) );
  BUFx3_ASAP7_75t_R register___U12664 ( .A(register__n9037), .Y(register__n8372) );
  BUFx4f_ASAP7_75t_R register___U12665 ( .A(register__n9800), .Y(register__n9053) );
  BUFx4f_ASAP7_75t_R register___U12666 ( .A(register__n9800), .Y(register__n9054) );
  BUFx2_ASAP7_75t_R register___U12667 ( .A(Reg_data[772]), .Y(register__n8373) );
  BUFx2_ASAP7_75t_R register___U12668 ( .A(Reg_data[281]), .Y(register__net98859) );
  BUFx2_ASAP7_75t_R register___U12669 ( .A(Reg_data[107]), .Y(register__net98847) );
  BUFx6f_ASAP7_75t_R register___U12670 ( .A(register__net89673), .Y(register__net98851) );
  BUFx4f_ASAP7_75t_R register___U12671 ( .A(register__net104013), .Y(register__net89673) );
  BUFx2_ASAP7_75t_R register___U12672 ( .A(Reg_data[126]), .Y(register__n8374) );
  BUFx4f_ASAP7_75t_R register___U12673 ( .A(register__n8377), .Y(register__n8375) );
  BUFx6f_ASAP7_75t_R register___U12674 ( .A(register__n8378), .Y(register__n8376) );
  BUFx3_ASAP7_75t_R register___U12675 ( .A(register__n10138), .Y(register__n8377) );
  BUFx6f_ASAP7_75t_R register___U12676 ( .A(register__n10138), .Y(register__n8378) );
  BUFx6f_ASAP7_75t_R register___U12677 ( .A(register__n10139), .Y(register__n10138) );
  BUFx4f_ASAP7_75t_R register___U12678 ( .A(register__n8021), .Y(register__n10139) );
  BUFx2_ASAP7_75t_R register___U12679 ( .A(Reg_data[556]), .Y(register__n8379) );
  BUFx2_ASAP7_75t_R register___U12680 ( .A(Reg_data[839]), .Y(register__net98827) );
  BUFx2_ASAP7_75t_R register___U12681 ( .A(Reg_data[279]), .Y(register__n8380) );
  INVx1_ASAP7_75t_R register___U12682 ( .A(register__n7348), .Y(register__n8381) );
  INVx1_ASAP7_75t_R register___U12683 ( .A(register__n7112), .Y(register__n8383) );
  BUFx3_ASAP7_75t_R register___U12684 ( .A(register__n8385), .Y(register__n8384) );
  BUFx2_ASAP7_75t_R register___U12685 ( .A(Reg_data[931]), .Y(register__n8385) );
  BUFx3_ASAP7_75t_R register___U12686 ( .A(register__net98690), .Y(register__net98689) );
  BUFx2_ASAP7_75t_R register___U12687 ( .A(Reg_data[914]), .Y(register__net98690) );
  BUFx3_ASAP7_75t_R register___U12688 ( .A(register__n8387), .Y(register__n8386) );
  BUFx2_ASAP7_75t_R register___U12689 ( .A(Reg_data[896]), .Y(register__n8387) );
  BUFx3_ASAP7_75t_R register___U12690 ( .A(register__n8389), .Y(register__n8388) );
  BUFx2_ASAP7_75t_R register___U12691 ( .A(Reg_data[854]), .Y(register__n8389) );
  BUFx3_ASAP7_75t_R register___U12692 ( .A(register__net98678), .Y(register__net98677) );
  BUFx2_ASAP7_75t_R register___U12693 ( .A(Reg_data[838]), .Y(register__net98678) );
  BUFx3_ASAP7_75t_R register___U12694 ( .A(register__net98674), .Y(register__net98673) );
  BUFx2_ASAP7_75t_R register___U12695 ( .A(Reg_data[837]), .Y(register__net98674) );
  BUFx3_ASAP7_75t_R register___U12696 ( .A(register__n8391), .Y(register__n8390) );
  BUFx2_ASAP7_75t_R register___U12697 ( .A(Reg_data[834]), .Y(register__n8391) );
  BUFx3_ASAP7_75t_R register___U12698 ( .A(register__n8393), .Y(register__n8392) );
  BUFx2_ASAP7_75t_R register___U12699 ( .A(Reg_data[789]), .Y(register__n8393) );
  BUFx3_ASAP7_75t_R register___U12700 ( .A(register__n8395), .Y(register__n8394) );
  BUFx2_ASAP7_75t_R register___U12701 ( .A(Reg_data[786]), .Y(register__n8395) );
  BUFx3_ASAP7_75t_R register___U12702 ( .A(register__net98658), .Y(register__net98657) );
  BUFx2_ASAP7_75t_R register___U12703 ( .A(Reg_data[774]), .Y(register__net98658) );
  BUFx3_ASAP7_75t_R register___U12704 ( .A(register__n8397), .Y(register__n8396) );
  BUFx2_ASAP7_75t_R register___U12705 ( .A(Reg_data[770]), .Y(register__n8397) );
  BUFx3_ASAP7_75t_R register___U12706 ( .A(register__n8399), .Y(register__n8398) );
  BUFx2_ASAP7_75t_R register___U12707 ( .A(Reg_data[768]), .Y(register__n8399) );
  BUFx3_ASAP7_75t_R register___U12708 ( .A(register__n8401), .Y(register__n8400) );
  BUFx2_ASAP7_75t_R register___U12709 ( .A(Reg_data[643]), .Y(register__n8401) );
  BUFx3_ASAP7_75t_R register___U12710 ( .A(register__n8403), .Y(register__n8402) );
  BUFx2_ASAP7_75t_R register___U12711 ( .A(Reg_data[597]), .Y(register__n8403) );
  BUFx3_ASAP7_75t_R register___U12712 ( .A(register__net98638), .Y(register__net98637) );
  BUFx2_ASAP7_75t_R register___U12713 ( .A(Reg_data[582]), .Y(register__net98638) );
  BUFx3_ASAP7_75t_R register___U12714 ( .A(register__net98634), .Y(register__net98633) );
  BUFx2_ASAP7_75t_R register___U12715 ( .A(Reg_data[409]), .Y(register__net98634) );
  BUFx3_ASAP7_75t_R register___U12716 ( .A(register__n8405), .Y(register__n8404) );
  BUFx2_ASAP7_75t_R register___U12717 ( .A(Reg_data[404]), .Y(register__n8405) );
  BUFx3_ASAP7_75t_R register___U12718 ( .A(register__n8407), .Y(register__n8406) );
  BUFx2_ASAP7_75t_R register___U12719 ( .A(Reg_data[322]), .Y(register__n8407) );
  BUFx3_ASAP7_75t_R register___U12720 ( .A(register__net98622), .Y(register__net98621) );
  BUFx2_ASAP7_75t_R register___U12721 ( .A(Reg_data[313]), .Y(register__net98622) );
  BUFx3_ASAP7_75t_R register___U12722 ( .A(register__n8409), .Y(register__n8408) );
  BUFx2_ASAP7_75t_R register___U12723 ( .A(Reg_data[308]), .Y(register__n8409) );
  BUFx3_ASAP7_75t_R register___U12724 ( .A(register__n8411), .Y(register__n8410) );
  BUFx2_ASAP7_75t_R register___U12725 ( .A(Reg_data[274]), .Y(register__n8411) );
  BUFx3_ASAP7_75t_R register___U12726 ( .A(register__n8413), .Y(register__n8412) );
  BUFx2_ASAP7_75t_R register___U12727 ( .A(Reg_data[256]), .Y(register__n8413) );
  BUFx3_ASAP7_75t_R register___U12728 ( .A(register__n8415), .Y(register__n8414) );
  BUFx2_ASAP7_75t_R register___U12729 ( .A(Reg_data[168]), .Y(register__n8415) );
  BUFx12f_ASAP7_75t_R register___U12730 ( .A(register__n7370), .Y(register__n8416) );
  BUFx12f_ASAP7_75t_R register___U12731 ( .A(register__n8416), .Y(register__n10008) );
  BUFx3_ASAP7_75t_R register___U12732 ( .A(register__net98599), .Y(register__net98598) );
  BUFx2_ASAP7_75t_R register___U12733 ( .A(Reg_data[166]), .Y(register__net98599) );
  BUFx3_ASAP7_75t_R register___U12734 ( .A(register__n8418), .Y(register__n8417) );
  BUFx2_ASAP7_75t_R register___U12735 ( .A(Reg_data[86]), .Y(register__n8418) );
  BUFx3_ASAP7_75t_R register___U12736 ( .A(register__n8420), .Y(register__n8419) );
  BUFx2_ASAP7_75t_R register___U12737 ( .A(Reg_data[85]), .Y(register__n8420) );
  BUFx3_ASAP7_75t_R register___U12738 ( .A(register__n8422), .Y(register__n8421) );
  BUFx2_ASAP7_75t_R register___U12739 ( .A(Reg_data[82]), .Y(register__n8422) );
  BUFx3_ASAP7_75t_R register___U12740 ( .A(register__net98583), .Y(register__net98582) );
  BUFx2_ASAP7_75t_R register___U12741 ( .A(Reg_data[70]), .Y(register__net98583) );
  BUFx3_ASAP7_75t_R register___U12742 ( .A(register__net98579), .Y(register__net98578) );
  BUFx2_ASAP7_75t_R register___U12743 ( .A(Reg_data[69]), .Y(register__net98579) );
  BUFx3_ASAP7_75t_R register___U12744 ( .A(register__n8424), .Y(register__n8423) );
  BUFx2_ASAP7_75t_R register___U12745 ( .A(Reg_data[66]), .Y(register__n8424) );
  BUFx3_ASAP7_75t_R register___U12746 ( .A(register__n8426), .Y(register__n8425) );
  BUFx2_ASAP7_75t_R register___U12747 ( .A(Reg_data[64]), .Y(register__n8426) );
  BUFx3_ASAP7_75t_R register___U12748 ( .A(register__n8428), .Y(register__n8427) );
  BUFx2_ASAP7_75t_R register___U12749 ( .A(Reg_data[872]), .Y(register__n8428) );
  BUFx3_ASAP7_75t_R register___U12750 ( .A(register__n8430), .Y(register__n8429) );
  BUFx2_ASAP7_75t_R register___U12751 ( .A(Reg_data[2]), .Y(register__n8430) );
  BUFx3_ASAP7_75t_R register___U12752 ( .A(register__n8432), .Y(register__n8431) );
  BUFx2_ASAP7_75t_R register___U12753 ( .A(Reg_data[0]), .Y(register__n8432) );
  BUFx3_ASAP7_75t_R register___U12754 ( .A(register__net98554), .Y(register__net98553) );
  BUFx2_ASAP7_75t_R register___U12755 ( .A(Reg_data[217]), .Y(register__net98554) );
  BUFx3_ASAP7_75t_R register___U12756 ( .A(register__n8434), .Y(register__n8433) );
  BUFx2_ASAP7_75t_R register___U12757 ( .A(Reg_data[21]), .Y(register__n8434) );
  BUFx3_ASAP7_75t_R register___U12758 ( .A(register__net98543), .Y(register__net98542) );
  BUFx2_ASAP7_75t_R register___U12759 ( .A(Reg_data[57]), .Y(register__net98543) );
  BUFx12f_ASAP7_75t_R register___U12760 ( .A(register__net89742), .Y(register__net89741) );
  BUFx3_ASAP7_75t_R register___U12761 ( .A(register__n8436), .Y(register__n8435) );
  BUFx2_ASAP7_75t_R register___U12762 ( .A(Reg_data[208]), .Y(register__n8436) );
  BUFx3_ASAP7_75t_R register___U12763 ( .A(register__n8438), .Y(register__n8437) );
  BUFx2_ASAP7_75t_R register___U12764 ( .A(Reg_data[194]), .Y(register__n8438) );
  BUFx3_ASAP7_75t_R register___U12765 ( .A(register__net98531), .Y(register__net98530) );
  BUFx2_ASAP7_75t_R register___U12766 ( .A(Reg_data[779]), .Y(register__net98531) );
  BUFx3_ASAP7_75t_R register___U12767 ( .A(register__net98527), .Y(register__net98526) );
  BUFx2_ASAP7_75t_R register___U12768 ( .A(Reg_data[75]), .Y(register__net98527) );
  BUFx3_ASAP7_75t_R register___U12769 ( .A(register__n8440), .Y(register__n8439) );
  BUFx2_ASAP7_75t_R register___U12770 ( .A(Reg_data[969]), .Y(register__n8440) );
  BUFx3_ASAP7_75t_R register___U12771 ( .A(register__net98519), .Y(register__net98518) );
  BUFx2_ASAP7_75t_R register___U12772 ( .A(Reg_data[600]), .Y(register__net98519) );
  BUFx3_ASAP7_75t_R register___U12773 ( .A(register__net98509), .Y(register__net98508) );
  BUFx2_ASAP7_75t_R register___U12774 ( .A(Reg_data[651]), .Y(register__net98509) );
  BUFx4f_ASAP7_75t_R register___U12775 ( .A(register__net89601), .Y(register__net98510) );
  BUFx2_ASAP7_75t_R register___U12776 ( .A(register__net89601), .Y(register__net98512) );
  BUFx4f_ASAP7_75t_R register___U12777 ( .A(register__net104011), .Y(register__net98498) );
  BUFx2_ASAP7_75t_R register___U12778 ( .A(Reg_data[88]), .Y(register__net98499) );
  BUFx12f_ASAP7_75t_R register___U12779 ( .A(register__net98501), .Y(register__net91331) );
  BUFx12f_ASAP7_75t_R register___U12780 ( .A(register__net91332), .Y(register__net98501) );
  BUFx6f_ASAP7_75t_R register___U12781 ( .A(register__net98498), .Y(register__net91332) );
  BUFx3_ASAP7_75t_R register___U12782 ( .A(register__net98495), .Y(register__net98494) );
  BUFx2_ASAP7_75t_R register___U12783 ( .A(Reg_data[335]), .Y(register__net98495) );
  BUFx3_ASAP7_75t_R register___U12784 ( .A(register__n8442), .Y(register__n8441) );
  BUFx2_ASAP7_75t_R register___U12785 ( .A(Reg_data[588]), .Y(register__n8442) );
  BUFx3_ASAP7_75t_R register___U12786 ( .A(register__n8444), .Y(register__n8443) );
  BUFx2_ASAP7_75t_R register___U12787 ( .A(Reg_data[795]), .Y(register__n8444) );
  BUFx3_ASAP7_75t_R register___U12788 ( .A(register__n8446), .Y(register__n8445) );
  BUFx2_ASAP7_75t_R register___U12789 ( .A(Reg_data[557]), .Y(register__n8446) );
  BUFx12f_ASAP7_75t_R register___U12790 ( .A(register__n10133), .Y(register__n8447) );
  BUFx12f_ASAP7_75t_R register___U12791 ( .A(register__n8447), .Y(register__n10132) );
  BUFx3_ASAP7_75t_R register___U12792 ( .A(register__n8449), .Y(register__n8448) );
  BUFx2_ASAP7_75t_R register___U12793 ( .A(Reg_data[30]), .Y(register__n8449) );
  BUFx3_ASAP7_75t_R register___U12794 ( .A(register__n8451), .Y(register__n8450) );
  BUFx2_ASAP7_75t_R register___U12795 ( .A(Reg_data[14]), .Y(register__n8451) );
  BUFx3_ASAP7_75t_R register___U12796 ( .A(register__n8453), .Y(register__n8452) );
  BUFx2_ASAP7_75t_R register___U12797 ( .A(Reg_data[653]), .Y(register__n8453) );
  BUFx4f_ASAP7_75t_R register___U12798 ( .A(register__n10150), .Y(register__n8454) );
  BUFx2_ASAP7_75t_R register___U12799 ( .A(register__n10150), .Y(register__n8455) );
  BUFx2_ASAP7_75t_R register___U12800 ( .A(register__n10150), .Y(register__n8456) );
  BUFx2_ASAP7_75t_R register___U12801 ( .A(Reg_data[481]), .Y(register__n8458) );
  BUFx3_ASAP7_75t_R register___U12802 ( .A(register__n8460), .Y(register__n8459) );
  BUFx2_ASAP7_75t_R register___U12803 ( .A(Reg_data[844]), .Y(register__n8460) );
  BUFx3_ASAP7_75t_R register___U12804 ( .A(register__n8462), .Y(register__n8461) );
  BUFx2_ASAP7_75t_R register___U12805 ( .A(Reg_data[204]), .Y(register__n8462) );
  BUFx3_ASAP7_75t_R register___U12806 ( .A(register__n8464), .Y(register__n8463) );
  BUFx2_ASAP7_75t_R register___U12807 ( .A(Reg_data[12]), .Y(register__n8464) );
  BUFx3_ASAP7_75t_R register___U12808 ( .A(register__n8466), .Y(register__n8465) );
  BUFx2_ASAP7_75t_R register___U12809 ( .A(Reg_data[94]), .Y(register__n8466) );
  BUFx3_ASAP7_75t_R register___U12810 ( .A(register__n8468), .Y(register__n8467) );
  BUFx2_ASAP7_75t_R register___U12811 ( .A(Reg_data[78]), .Y(register__n8468) );
  BUFx3_ASAP7_75t_R register___U12812 ( .A(register__n8470), .Y(register__n8469) );
  BUFx2_ASAP7_75t_R register___U12813 ( .A(Reg_data[350]), .Y(register__n8470) );
  BUFx4f_ASAP7_75t_R register___U12814 ( .A(register__net108335), .Y(register__net98422) );
  BUFx2_ASAP7_75t_R register___U12815 ( .A(Reg_data[472]), .Y(register__net98423) );
  BUFx12f_ASAP7_75t_R register___U12816 ( .A(register__net90538), .Y(register__net90537) );
  BUFx6f_ASAP7_75t_R register___U12817 ( .A(register__net98422), .Y(register__net90538) );
  BUFx3_ASAP7_75t_R register___U12818 ( .A(register__net98416), .Y(register__net98415) );
  BUFx2_ASAP7_75t_R register___U12819 ( .A(Reg_data[440]), .Y(register__net98416) );
  BUFx12f_ASAP7_75t_R register___U12820 ( .A(register__net88417), .Y(register__net88416) );
  BUFx4f_ASAP7_75t_R register___U12821 ( .A(register__net108333), .Y(register__net98407) );
  BUFx2_ASAP7_75t_R register___U12822 ( .A(Reg_data[943]), .Y(register__net98408) );
  BUFx12f_ASAP7_75t_R register___U12823 ( .A(register__net90530), .Y(register__net90529) );
  BUFx6f_ASAP7_75t_R register___U12824 ( .A(register__net98407), .Y(register__net90530) );
  BUFx3_ASAP7_75t_R register___U12825 ( .A(register__net98401), .Y(register__net98400) );
  BUFx2_ASAP7_75t_R register___U12826 ( .A(Reg_data[175]), .Y(register__net98401) );
  BUFx12f_ASAP7_75t_R register___U12827 ( .A(register__net89406), .Y(register__net89405) );
  BUFx3_ASAP7_75t_R register___U12828 ( .A(register__net98397), .Y(register__net98396) );
  BUFx2_ASAP7_75t_R register___U12829 ( .A(Reg_data[463]), .Y(register__net98397) );
  BUFx3_ASAP7_75t_R register___U12830 ( .A(register__n8472), .Y(register__n8471) );
  BUFx2_ASAP7_75t_R register___U12831 ( .A(Reg_data[483]), .Y(register__n8472) );
  BUFx3_ASAP7_75t_R register___U12832 ( .A(register__n8474), .Y(register__n8473) );
  BUFx2_ASAP7_75t_R register___U12833 ( .A(Reg_data[571]), .Y(register__n8474) );
  BUFx4f_ASAP7_75t_R register___U12834 ( .A(register__n8022), .Y(register__n8475) );
  BUFx2_ASAP7_75t_R register___U12835 ( .A(Reg_data[679]), .Y(register__n8476) );
  BUFx12f_ASAP7_75t_R register___U12836 ( .A(register__n10188), .Y(register__n8477) );
  BUFx12f_ASAP7_75t_R register___U12837 ( .A(register__n8477), .Y(register__n10187) );
  BUFx6f_ASAP7_75t_R register___U12838 ( .A(register__n8475), .Y(register__n10188) );
  BUFx3_ASAP7_75t_R register___U12839 ( .A(register__n8479), .Y(register__n8478) );
  BUFx2_ASAP7_75t_R register___U12840 ( .A(Reg_data[455]), .Y(register__n8479) );
  BUFx12f_ASAP7_75t_R register___U12841 ( .A(register__n9787), .Y(register__n8480) );
  BUFx12f_ASAP7_75t_R register___U12842 ( .A(register__n8480), .Y(register__n9786) );
  BUFx3_ASAP7_75t_R register___U12843 ( .A(register__n8482), .Y(register__n8481) );
  BUFx2_ASAP7_75t_R register___U12844 ( .A(Reg_data[487]), .Y(register__n8482) );
  BUFx12f_ASAP7_75t_R register___U12845 ( .A(register__n9298), .Y(register__n8483) );
  BUFx12f_ASAP7_75t_R register___U12846 ( .A(register__n8483), .Y(register__n9297) );
  BUFx4f_ASAP7_75t_R register___U12847 ( .A(register__n5176), .Y(register__n8484) );
  BUFx2_ASAP7_75t_R register___U12848 ( .A(Reg_data[958]), .Y(register__n8485) );
  BUFx12f_ASAP7_75t_R register___U12849 ( .A(register__n9805), .Y(register__n9804) );
  BUFx6f_ASAP7_75t_R register___U12850 ( .A(register__n8484), .Y(register__n9805) );
  BUFx3_ASAP7_75t_R register___U12851 ( .A(register__n8487), .Y(register__n8486) );
  BUFx2_ASAP7_75t_R register___U12852 ( .A(Reg_data[190]), .Y(register__n8487) );
  BUFx12f_ASAP7_75t_R register___U12853 ( .A(register__n7378), .Y(register__n10203) );
  BUFx3_ASAP7_75t_R register___U12854 ( .A(register__n8489), .Y(register__n8488) );
  BUFx2_ASAP7_75t_R register___U12855 ( .A(Reg_data[718]), .Y(register__n8489) );
  BUFx4f_ASAP7_75t_R register___U12856 ( .A(register__n10221), .Y(register__n8490) );
  BUFx2_ASAP7_75t_R register___U12857 ( .A(register__n10221), .Y(register__n8491) );
  BUFx3_ASAP7_75t_R register___U12858 ( .A(register__n8494), .Y(register__n8493) );
  BUFx2_ASAP7_75t_R register___U12859 ( .A(Reg_data[798]), .Y(register__n8494) );
  BUFx4f_ASAP7_75t_R register___U12860 ( .A(register__n8023), .Y(register__n8495) );
  BUFx2_ASAP7_75t_R register___U12861 ( .A(Reg_data[862]), .Y(register__n8496) );
  BUFx12f_ASAP7_75t_R register___U12862 ( .A(register__n8498), .Y(register__n8497) );
  BUFx12f_ASAP7_75t_R register___U12863 ( .A(register__n10390), .Y(register__n8498) );
  BUFx12f_ASAP7_75t_R register___U12864 ( .A(register__n8497), .Y(register__n10389) );
  BUFx6f_ASAP7_75t_R register___U12865 ( .A(register__n8495), .Y(register__n10390) );
  BUFx3_ASAP7_75t_R register___U12866 ( .A(register__n8500), .Y(register__n8499) );
  BUFx2_ASAP7_75t_R register___U12867 ( .A(Reg_data[716]), .Y(register__n8500) );
  BUFx12f_ASAP7_75t_R register___U12868 ( .A(register__n10234), .Y(register__n8501) );
  BUFx12f_ASAP7_75t_R register___U12869 ( .A(register__n8501), .Y(register__n10233) );
  BUFx3_ASAP7_75t_R register___U12870 ( .A(register__n8503), .Y(register__n8502) );
  BUFx2_ASAP7_75t_R register___U12871 ( .A(Reg_data[659]), .Y(register__n8503) );
  BUFx4f_ASAP7_75t_R register___U12872 ( .A(register__n10247), .Y(register__n8504) );
  BUFx2_ASAP7_75t_R register___U12873 ( .A(register__n10247), .Y(register__n8505) );
  BUFx2_ASAP7_75t_R register___U12874 ( .A(register__n10247), .Y(register__n8506) );
  BUFx3_ASAP7_75t_R register___U12875 ( .A(register__net98311), .Y(register__net98310) );
  BUFx2_ASAP7_75t_R register___U12876 ( .A(Reg_data[859]), .Y(register__net98311) );
  BUFx3_ASAP7_75t_R register___U12877 ( .A(register__n8508), .Y(register__n8507) );
  BUFx2_ASAP7_75t_R register___U12878 ( .A(Reg_data[215]), .Y(register__n8508) );
  BUFx3_ASAP7_75t_R register___U12879 ( .A(register__n10269), .Y(register__n8509) );
  BUFx2_ASAP7_75t_R register___U12880 ( .A(register__n10269), .Y(register__n8510) );
  BUFx4f_ASAP7_75t_R register___U12881 ( .A(register__n10269), .Y(register__n8511) );
  BUFx3_ASAP7_75t_R register___U12882 ( .A(register__n8513), .Y(register__n8512) );
  BUFx2_ASAP7_75t_R register___U12883 ( .A(Reg_data[922]), .Y(register__n8513) );
  BUFx2_ASAP7_75t_R register___U12884 ( .A(register__n9309), .Y(register__n8514) );
  BUFx2_ASAP7_75t_R register___U12885 ( .A(register__n9309), .Y(register__n8515) );
  BUFx4f_ASAP7_75t_R register___U12886 ( .A(register__n9309), .Y(register__n8516) );
  BUFx3_ASAP7_75t_R register___U12887 ( .A(register__n8518), .Y(register__n8517) );
  BUFx2_ASAP7_75t_R register___U12888 ( .A(Reg_data[191]), .Y(register__n8518) );
  BUFx12f_ASAP7_75t_R register___U12889 ( .A(register__n10296), .Y(register__n8519) );
  BUFx12f_ASAP7_75t_R register___U12890 ( .A(register__n8519), .Y(register__n10295) );
  BUFx3_ASAP7_75t_R register___U12891 ( .A(register__n8521), .Y(register__n8520) );
  BUFx2_ASAP7_75t_R register___U12892 ( .A(Reg_data[713]), .Y(register__n8521) );
  BUFx4f_ASAP7_75t_R register___U12893 ( .A(register__n10299), .Y(register__n8522) );
  BUFx2_ASAP7_75t_R register___U12894 ( .A(register__n10299), .Y(register__n8523) );
  BUFx3_ASAP7_75t_R register___U12895 ( .A(register__n8526), .Y(register__n8525) );
  BUFx2_ASAP7_75t_R register___U12896 ( .A(Reg_data[396]), .Y(register__n8526) );
  BUFx2_ASAP7_75t_R register___U12897 ( .A(register__n9877), .Y(register__n8527) );
  BUFx2_ASAP7_75t_R register___U12898 ( .A(register__n9877), .Y(register__n8528) );
  BUFx4f_ASAP7_75t_R register___U12899 ( .A(register__n9877), .Y(register__n8529) );
  BUFx3_ASAP7_75t_R register___U12900 ( .A(register__n8531), .Y(register__n8530) );
  BUFx2_ASAP7_75t_R register___U12901 ( .A(Reg_data[428]), .Y(register__n8531) );
  BUFx12f_ASAP7_75t_R register___U12902 ( .A(register__n9880), .Y(register__n8532) );
  BUFx12f_ASAP7_75t_R register___U12903 ( .A(register__n8532), .Y(register__n9879) );
  BUFx4f_ASAP7_75t_R register___U12904 ( .A(register__n6280), .Y(register__n8533) );
  BUFx2_ASAP7_75t_R register___U12905 ( .A(Reg_data[657]), .Y(register__n8534) );
  BUFx12f_ASAP7_75t_R register___U12906 ( .A(register__n10314), .Y(register__n8535) );
  BUFx12f_ASAP7_75t_R register___U12907 ( .A(register__n8535), .Y(register__n10313) );
  BUFx6f_ASAP7_75t_R register___U12908 ( .A(register__n8533), .Y(register__n10314) );
  BUFx3_ASAP7_75t_R register___U12909 ( .A(register__n8537), .Y(register__n8536) );
  BUFx2_ASAP7_75t_R register___U12910 ( .A(Reg_data[401]), .Y(register__n8537) );
  BUFx2_ASAP7_75t_R register___U12911 ( .A(register__n9885), .Y(register__n8538) );
  BUFx2_ASAP7_75t_R register___U12912 ( .A(register__n9885), .Y(register__n8539) );
  BUFx4f_ASAP7_75t_R register___U12913 ( .A(register__n9885), .Y(register__n8540) );
  BUFx3_ASAP7_75t_R register___U12914 ( .A(register__n8542), .Y(register__n8541) );
  BUFx2_ASAP7_75t_R register___U12915 ( .A(Reg_data[465]), .Y(register__n8542) );
  BUFx12f_ASAP7_75t_R register___U12916 ( .A(register__n9890), .Y(register__n8543) );
  BUFx12f_ASAP7_75t_R register___U12917 ( .A(register__n8543), .Y(register__n9889) );
  BUFx3_ASAP7_75t_R register___U12918 ( .A(register__net98225), .Y(register__net98224) );
  BUFx2_ASAP7_75t_R register___U12919 ( .A(Reg_data[664]), .Y(register__net98225) );
  BUFx4f_ASAP7_75t_R register___U12920 ( .A(register__net103999), .Y(register__net98214) );
  BUFx2_ASAP7_75t_R register___U12921 ( .A(Reg_data[856]), .Y(register__net98215) );
  BUFx12f_ASAP7_75t_R register___U12922 ( .A(register__net98217), .Y(register__net88785) );
  BUFx12f_ASAP7_75t_R register___U12923 ( .A(register__net88786), .Y(register__net98217) );
  BUFx6f_ASAP7_75t_R register___U12924 ( .A(register__net98214), .Y(register__net88786) );
  BUFx3_ASAP7_75t_R register___U12925 ( .A(register__net98211), .Y(register__net98210) );
  BUFx2_ASAP7_75t_R register___U12926 ( .A(Reg_data[765]), .Y(register__net98211) );
  BUFx3_ASAP7_75t_R register___U12927 ( .A(register__net98207), .Y(register__net98206) );
  BUFx2_ASAP7_75t_R register___U12928 ( .A(Reg_data[925]), .Y(register__net98207) );
  BUFx3_ASAP7_75t_R register___U12929 ( .A(register__net98202), .Y(register__net98201) );
  BUFx2_ASAP7_75t_R register___U12930 ( .A(Reg_data[957]), .Y(register__net98202) );
  BUFx3_ASAP7_75t_R register___U12931 ( .A(register__net98192), .Y(register__net98191) );
  BUFx2_ASAP7_75t_R register___U12932 ( .A(Reg_data[541]), .Y(register__net98192) );
  BUFx4f_ASAP7_75t_R register___U12933 ( .A(register__net89017), .Y(register__net98193) );
  BUFx3_ASAP7_75t_R register___U12934 ( .A(register__net98185), .Y(register__net98184) );
  BUFx2_ASAP7_75t_R register___U12935 ( .A(Reg_data[701]), .Y(register__net98185) );
  BUFx12f_ASAP7_75t_R register___U12936 ( .A(register__net89002), .Y(register__net89001) );
  BUFx4f_ASAP7_75t_R register___U12937 ( .A(register__n3252), .Y(register__n8544) );
  BUFx2_ASAP7_75t_R register___U12938 ( .A(Reg_data[956]), .Y(register__n8545) );
  BUFx6f_ASAP7_75t_R register___U12939 ( .A(register__n8544), .Y(register__n9902) );
  BUFx3_ASAP7_75t_R register___U12940 ( .A(register__n8547), .Y(register__n8546) );
  BUFx2_ASAP7_75t_R register___U12941 ( .A(Reg_data[156]), .Y(register__n8547) );
  BUFx4f_ASAP7_75t_R register___U12942 ( .A(register__n10331), .Y(register__n8548) );
  BUFx2_ASAP7_75t_R register___U12943 ( .A(register__n10331), .Y(register__n8549) );
  BUFx3_ASAP7_75t_R register___U12944 ( .A(register__n10331), .Y(register__n8550) );
  BUFx3_ASAP7_75t_R register___U12945 ( .A(register__n8552), .Y(register__n8551) );
  BUFx2_ASAP7_75t_R register___U12946 ( .A(Reg_data[188]), .Y(register__n8552) );
  BUFx12f_ASAP7_75t_R register___U12947 ( .A(register__n5180), .Y(register__n10333) );
  BUFx3_ASAP7_75t_R register___U12948 ( .A(register__n8554), .Y(register__n8553) );
  BUFx2_ASAP7_75t_R register___U12949 ( .A(Reg_data[462]), .Y(register__n8554) );
  INVx2_ASAP7_75t_R register___U12950 ( .A(register__net94176), .Y(register__net98142) );
  BUFx6f_ASAP7_75t_R register___U12951 ( .A(register__net94177), .Y(register__net94176) );
  OA22x2_ASAP7_75t_R register___U12952 ( .A1(register__n12229), .A2(register__n1092), .B1(register__n9883), .B2(register__n11761), 
        .Y(register__n13074) );
  INVx1_ASAP7_75t_R register___U12953 ( .A(register__n4675), .Y(register__n8555) );
  OA22x2_ASAP7_75t_R register___U12954 ( .A1(register__net62656), .A2(register__n1755), .B1(register__n9891), .B2(register__n3334), .Y(register__n13116) );
  OA22x2_ASAP7_75t_R register___U12955 ( .A1(register__n12460), .A2(register__n1946), .B1(register__n6932), .B2(register__n1992), 
        .Y(register__n12801) );
  INVx4_ASAP7_75t_R register___U12956 ( .A(register__n12475), .Y(register__n12460) );
  INVx1_ASAP7_75t_R register___U12957 ( .A(register__n11027), .Y(register__n8557) );
  INVx1_ASAP7_75t_R register___U12958 ( .A(register__n4708), .Y(register__n8558) );
  BUFx12f_ASAP7_75t_R register___U12959 ( .A(register__n12076), .Y(register__n8563) );
  INVx1_ASAP7_75t_R register___U12960 ( .A(register__n5015), .Y(register__n8566) );
  INVx1_ASAP7_75t_R register___U12961 ( .A(register__n5017), .Y(register__n8567) );
  INVx1_ASAP7_75t_R register___U12962 ( .A(register__n5019), .Y(register__n8568) );
  INVx1_ASAP7_75t_R register___U12963 ( .A(register__n5261), .Y(register__n8570) );
  INVx1_ASAP7_75t_R register___U12964 ( .A(register__n5064), .Y(register__n8572) );
  INVx1_ASAP7_75t_R register___U12965 ( .A(register__n4228), .Y(register__n8573) );
  INVx1_ASAP7_75t_R register___U12966 ( .A(register__n4862), .Y(register__n8576) );
  INVx1_ASAP7_75t_R register___U12967 ( .A(register__n5558), .Y(register__n8577) );
  INVx1_ASAP7_75t_R register___U12968 ( .A(register__n11573), .Y(register__n8579) );
  INVx1_ASAP7_75t_R register___U12969 ( .A(register__n4099), .Y(register__n8581) );
  OA22x2_ASAP7_75t_R register___U12970 ( .A1(register__n12461), .A2(register__n104), .B1(register__n9061), .B2(register__n1100), 
        .Y(register__n12747) );
  OA22x2_ASAP7_75t_R register___U12971 ( .A1(register__n12426), .A2(register__n951), .B1(register__n10505), .B2(register__n959), 
        .Y(register__n13012) );
  INVx1_ASAP7_75t_R register___U12972 ( .A(register__n3585), .Y(register__n8583) );
  INVx3_ASAP7_75t_R register___U12973 ( .A(register__n8014), .Y(register__n8588) );
  INVx3_ASAP7_75t_R register___U12974 ( .A(register__n11349), .Y(register__n8589) );
  INVx3_ASAP7_75t_R register___U12975 ( .A(register__n10740), .Y(register__n8590) );
  INVx3_ASAP7_75t_R register___U12976 ( .A(register__n11500), .Y(register__n8591) );
  OA22x2_ASAP7_75t_R register___U12977 ( .A1(register__n11928), .A2(register__n462), .B1(register__n9997), .B2(register__n463), 
        .Y(register__n12949) );
  INVx1_ASAP7_75t_R register___U12978 ( .A(register__n5753), .Y(register__n8592) );
  OA22x2_ASAP7_75t_R register___U12979 ( .A1(register__n11955), .A2(register__n891), .B1(register__n10495), .B2(register__n903), 
        .Y(register__n13063) );
  INVx1_ASAP7_75t_R register___U12980 ( .A(register__n5757), .Y(register__n8593) );
  OA22x2_ASAP7_75t_R register___U12981 ( .A1(register__n12087), .A2(register__n462), .B1(register__n10421), .B2(register__n474), 
        .Y(register__n12940) );
  OA22x2_ASAP7_75t_R register___U12982 ( .A1(register__net63006), .A2(register__n339), .B1(register__n9351), .B2(register__n68), 
        .Y(register__n12721) );
  OA22x2_ASAP7_75t_R register___U12983 ( .A1(register__net62666), .A2(register__n109), .B1(register__n9321), .B2(register__n5501), 
        .Y(register__n12831) );
  OA22x2_ASAP7_75t_R register___U12984 ( .A1(register__n12203), .A2(register__n182), .B1(register__n10481), .B2(register__n213), 
        .Y(register__n12676) );
  INVx1_ASAP7_75t_R register___U12985 ( .A(register__n12676), .Y(register__n8596) );
  OA22x2_ASAP7_75t_R register___U12986 ( .A1(register__n12346), .A2(register__n337), .B1(register__n10509), .B2(register__n342), 
        .Y(register__n12726) );
  OA22x2_ASAP7_75t_R register___U12987 ( .A1(register__n12202), .A2(register__n1794), .B1(register__n9355), .B2(register__n1625), 
        .Y(register__n12761) );
  OA22x2_ASAP7_75t_R register___U12988 ( .A1(register__n12458), .A2(register__n1973), .B1(register__n9417), .B2(register__n2136), 
        .Y(register__n12889) );
  OA22x2_ASAP7_75t_R register___U12989 ( .A1(register__net63006), .A2(register__n1643), .B1(register__n10473), .B2(
        n1638), .Y(register__n12750) );
  INVx1_ASAP7_75t_R register___U12990 ( .A(register__n12750), .Y(register__n8598) );
  OA22x2_ASAP7_75t_R register___U12991 ( .A1(register__n12233), .A2(register__n2220), .B1(register__n10315), .B2(register__n1463), 
        .Y(register__n12785) );
  OA22x2_ASAP7_75t_R register___U12992 ( .A1(register__net62658), .A2(register__n2144), .B1(register__n9217), .B2(register__n1207), .Y(register__n13088) );
  INVx1_ASAP7_75t_R register___U12993 ( .A(register__n4092), .Y(register__n8599) );
  OA22x2_ASAP7_75t_R register___U12994 ( .A1(register__n12028), .A2(register__n1098), .B1(register__n10444), .B2(register__n3508), 
        .Y(register__n12797) );
  OA22x2_ASAP7_75t_R register___U12995 ( .A1(register__n12257), .A2(register__n109), .B1(register__n9959), .B2(register__n5503), 
        .Y(register__n12842) );
  INVx1_ASAP7_75t_R register___U12996 ( .A(register__n7120), .Y(register__n8602) );
  OA22x2_ASAP7_75t_R register___U12997 ( .A1(register__net64766), .A2(register__n109), .B1(register__net90041), .B2(
        n5660), .Y(register__n12854) );
  OA22x2_ASAP7_75t_R register___U12998 ( .A1(register__n12027), .A2(register__n109), .B1(register__n9963), .B2(register__n12499), 
        .Y(register__n12857) );
  OA22x2_ASAP7_75t_R register___U12999 ( .A1(register__n11927), .A2(register__n1413), .B1(register__n9640), .B2(register__n1417), 
        .Y(register__n13009) );
  OA22x2_ASAP7_75t_R register___U13000 ( .A1(register__n12369), .A2(register__n951), .B1(register__n9642), .B2(register__n958), 
        .Y(register__n13018) );
  INVx1_ASAP7_75t_R register___U13001 ( .A(register__n4870), .Y(register__n8604) );
  OA22x2_ASAP7_75t_R register___U13002 ( .A1(register__n12341), .A2(register__n1092), .B1(register__n9670), .B2(register__n7336), 
        .Y(register__n13071) );
  BUFx12f_ASAP7_75t_R register___U13003 ( .A(register__n6523), .Y(register__n9674) );
  OA22x2_ASAP7_75t_R register___U13004 ( .A1(register__n11988), .A2(register__n1092), .B1(register__n9678), .B2(register__n7663), 
        .Y(register__n13086) );
  OA22x2_ASAP7_75t_R register___U13005 ( .A1(register__net63254), .A2(register__n109), .B1(register__net89649), .B2(
        n5502), .Y(register__n12837) );
  INVx1_ASAP7_75t_R register___U13006 ( .A(register__n4663), .Y(register__n8608) );
  OA22x2_ASAP7_75t_R register___U13007 ( .A1(register__n12086), .A2(register__n1414), .B1(register__n10432), .B2(register__n1418), 
        .Y(register__n13000) );
  OA22x2_ASAP7_75t_R register___U13008 ( .A1(register__n12234), .A2(register__n3719), .B1(register__n9543), .B2(register__n1163), 
        .Y(register__n13372) );
  OA22x2_ASAP7_75t_R register___U13009 ( .A1(register__net146308), .A2(register__n118), .B1(register__n9545), .B2(register__n1202), .Y(register__n13092) );
  INVx1_ASAP7_75t_R register___U13010 ( .A(register__n6791), .Y(register__n8610) );
  OA22x2_ASAP7_75t_R register___U13011 ( .A1(register__n12088), .A2(register__n109), .B1(register__n10167), .B2(register__n8358), 
        .Y(register__n12851) );
  OA22x2_ASAP7_75t_R register___U13012 ( .A1(register__n12091), .A2(register__n178), .B1(register__n7191), .B2(register__n207), 
        .Y(register__n12683) );
  INVx1_ASAP7_75t_R register___U13013 ( .A(register__n4671), .Y(register__n8611) );
  OA22x2_ASAP7_75t_R register___U13014 ( .A1(register__net63246), .A2(register__n1092), .B1(register__net90545), .B2(
        n11763), .Y(register__n13068) );
  INVx1_ASAP7_75t_R register___U13015 ( .A(register__n4881), .Y(register__n8612) );
  OA22x2_ASAP7_75t_R register___U13016 ( .A1(register__net64432), .A2(register__n2220), .B1(register__net93404), .B2(
        n485), .Y(register__n12790) );
  INVx3_ASAP7_75t_R register___U13017 ( .A(register__net64466), .Y(register__net64432) );
  OA22x2_ASAP7_75t_R register___U13018 ( .A1(register__n12084), .A2(register__n1092), .B1(register__n9849), .B2(register__n11757), 
        .Y(register__n13081) );
  INVx1_ASAP7_75t_R register___U13019 ( .A(register__n6799), .Y(register__n8613) );
  OA22x2_ASAP7_75t_R register___U13020 ( .A1(register__n12115), .A2(register__n1092), .B1(register__n8194), .B2(register__n6430), 
        .Y(register__n13079) );
  INVx1_ASAP7_75t_R register___U13021 ( .A(register__n4890), .Y(register__n8614) );
  OA22x2_ASAP7_75t_R register___U13022 ( .A1(register__net63258), .A2(register__n175), .B1(register__net90261), .B2(
        n213), .Y(register__n12668) );
  OA22x2_ASAP7_75t_R register___U13023 ( .A1(register__net63256), .A2(register__n2220), .B1(register__net89041), .B2(
        n11806), .Y(register__n12783) );
  OA22x2_ASAP7_75t_R register___U13024 ( .A1(register__n12430), .A2(register__n2220), .B1(register__n10337), .B2(register__n11807), .Y(register__n12779) );
  OA22x2_ASAP7_75t_R register___U13025 ( .A1(register__n12147), .A2(register__n1569), .B1(register__n10377), .B2(register__n1189), 
        .Y(register__n13102) );
  OA22x2_ASAP7_75t_R register___U13026 ( .A1(register__n12260), .A2(register__n194), .B1(register__n9613), .B2(register__n205), 
        .Y(register__n12674) );
  INVx1_ASAP7_75t_R register___U13027 ( .A(register__n4293), .Y(register__n8616) );
  OA22x2_ASAP7_75t_R register___U13028 ( .A1(register__net64856), .A2(register__n181), .B1(register__net90997), .B2(
        n205), .Y(register__n12686) );
  INVx1_ASAP7_75t_R register___U13029 ( .A(register__n12686), .Y(register__n8617) );
  OA22x2_ASAP7_75t_R register___U13030 ( .A1(register__n11960), .A2(register__n337), .B1(register__n6848), .B2(register__n345), 
        .Y(register__n12745) );
  INVx1_ASAP7_75t_R register___U13031 ( .A(register__n3577), .Y(register__n8618) );
  BUFx6f_ASAP7_75t_R register___U13032 ( .A(register__n12417), .Y(register__n12410) );
  BUFx6f_ASAP7_75t_R register___U13033 ( .A(register__n12415), .Y(register__n12408) );
  OA22x2_ASAP7_75t_R register___U13034 ( .A1(register__n12429), .A2(register__n109), .B1(register__n9367), .B2(register__n3307), 
        .Y(register__n12834) );
  OA22x2_ASAP7_75t_R register___U13035 ( .A1(register__n12458), .A2(register__n459), .B1(register__n10206), .B2(register__n471), 
        .Y(register__n12920) );
  INVx1_ASAP7_75t_R register___U13036 ( .A(register__n5783), .Y(register__n8621) );
  OA22x2_ASAP7_75t_R register___U13037 ( .A1(register__net62816), .A2(register__n1989), .B1(register__net91583), .B2(
        n11851), .Y(register__n13336) );
  OA22x2_ASAP7_75t_R register___U13038 ( .A1(register__net62836), .A2(register__n1946), .B1(register__net89005), .B2(
        n1992), .Y(register__n12802) );
  INVx1_ASAP7_75t_R register___U13039 ( .A(register__n12802), .Y(register__n8623) );
  OA22x2_ASAP7_75t_R register___U13040 ( .A1(register__n12431), .A2(register__n1647), .B1(register__n10475), .B2(register__n1627), 
        .Y(register__n12749) );
  OA22x2_ASAP7_75t_R register___U13041 ( .A1(register__n12457), .A2(register__n895), .B1(register__n9903), .B2(register__n907), 
        .Y(register__n13039) );
  INVx1_ASAP7_75t_R register___U13042 ( .A(register__n4619), .Y(register__n8628) );
  INVx1_ASAP7_75t_R register___U13043 ( .A(register__n4787), .Y(register__n8629) );
  INVx1_ASAP7_75t_R register___U13044 ( .A(register__n4789), .Y(register__n8630) );
  INVx1_ASAP7_75t_R register___U13045 ( .A(register__n4791), .Y(register__n8631) );
  INVx1_ASAP7_75t_R register___U13046 ( .A(register__n6516), .Y(register__n8632) );
  INVx1_ASAP7_75t_R register___U13047 ( .A(register__n6518), .Y(register__n8633) );
  INVx1_ASAP7_75t_R register___U13048 ( .A(register__n10902), .Y(register__n8634) );
  INVx1_ASAP7_75t_R register___U13049 ( .A(register__n5305), .Y(register__n8636) );
  INVx1_ASAP7_75t_R register___U13050 ( .A(register__n5397), .Y(register__n8637) );
  BUFx6f_ASAP7_75t_R register___U13051 ( .A(register__net127351), .Y(register__net64698) );
  BUFx6f_ASAP7_75t_R register___U13052 ( .A(register__net127351), .Y(register__net64704) );
  OA22x2_ASAP7_75t_R register___U13053 ( .A1(register__n12347), .A2(register__n185), .B1(register__n9609), .B2(register__n204), 
        .Y(register__n12671) );
  INVx1_ASAP7_75t_R register___U13054 ( .A(register__n5002), .Y(register__n8646) );
  OA22x2_ASAP7_75t_R register___U13055 ( .A1(register__n3501), .A2(register__n1415), .B1(register__n9638), .B2(register__n1417), 
        .Y(register__n13006) );
  INVx1_ASAP7_75t_R register___U13056 ( .A(register__n4134), .Y(register__n8647) );
  OA22x2_ASAP7_75t_R register___U13057 ( .A1(register__n12032), .A2(register__n1643), .B1(register__n9419), .B2(register__n1617), 
        .Y(register__n12773) );
  OA22x2_ASAP7_75t_R register___U13058 ( .A1(register__n12201), .A2(register__n1069), .B1(register__n9421), .B2(register__n81), 
        .Y(register__n12815) );
  INVx1_ASAP7_75t_R register___U13059 ( .A(register__n3611), .Y(register__n8649) );
  OA22x2_ASAP7_75t_R register___U13060 ( .A1(register__n12372), .A2(register__n1920), .B1(register__n9459), .B2(register__n1924), 
        .Y(register__n12867) );
  INVx1_ASAP7_75t_R register___U13061 ( .A(register__n5566), .Y(register__n8650) );
  OA22x2_ASAP7_75t_R register___U13062 ( .A1(register__n5351), .A2(register__n11885), .B1(register__n9463), .B2(register__n1952), 
        .Y(register__n12869) );
  INVx1_ASAP7_75t_R register___U13063 ( .A(register__n6238), .Y(register__n8651) );
  OA22x2_ASAP7_75t_R register___U13064 ( .A1(register__n12200), .A2(register__n2820), .B1(register__n9465), .B2(register__n1940), 
        .Y(register__n12873) );
  INVx1_ASAP7_75t_R register___U13065 ( .A(register__n4054), .Y(register__n8652) );
  OA22x2_ASAP7_75t_R register___U13066 ( .A1(register__n3644), .A2(register__n1923), .B1(register__n9469), .B2(register__n1937), 
        .Y(register__n12885) );
  INVx1_ASAP7_75t_R register___U13067 ( .A(register__n4056), .Y(register__n8653) );
  OA22x2_ASAP7_75t_R register___U13068 ( .A1(register__net142376), .A2(register__n892), .B1(register__net114453), .B2(
        n899), .Y(register__n13059) );
  OA22x2_ASAP7_75t_R register___U13069 ( .A1(register__n12315), .A2(register__n1565), .B1(register__n9471), .B2(register__n1210), 
        .Y(register__n13095) );
  OA22x2_ASAP7_75t_R register___U13070 ( .A1(register__net64758), .A2(register__n1567), .B1(register__net91447), .B2(
        n1185), .Y(register__n13109) );
  OA22x2_ASAP7_75t_R register___U13071 ( .A1(register__n11930), .A2(register__n118), .B1(register__n9473), .B2(register__n1203), 
        .Y(register__n13115) );
  OA22x2_ASAP7_75t_R register___U13072 ( .A1(register__n3467), .A2(register__n1140), .B1(register__n9475), .B2(register__n1058), 
        .Y(register__n13156) );
  INVx1_ASAP7_75t_R register___U13073 ( .A(register__n3738), .Y(register__n8656) );
  OA22x2_ASAP7_75t_R register___U13074 ( .A1(register__n12340), .A2(register__n1140), .B1(register__n9477), .B2(register__n1147), 
        .Y(register__n13157) );
  INVx1_ASAP7_75t_R register___U13075 ( .A(register__n3824), .Y(register__n8657) );
  OA22x2_ASAP7_75t_R register___U13076 ( .A1(register__net64352), .A2(register__n2822), .B1(register__net91347), .B2(
        n1930), .Y(register__n12877) );
  OA22x2_ASAP7_75t_R register___U13077 ( .A1(register__n12232), .A2(register__n109), .B1(register__n7142), .B2(register__n11800), 
        .Y(register__n12843) );
  INVx1_ASAP7_75t_R register___U13078 ( .A(register__n4665), .Y(register__n8659) );
  OA22x2_ASAP7_75t_R register___U13079 ( .A1(register__net64012), .A2(register__n665), .B1(register__net88628), .B2(register__n81), .Y(register__n12816) );
  BUFx12f_ASAP7_75t_R register___U13080 ( .A(register__n7779), .Y(register__n9527) );
  OA22x2_ASAP7_75t_R register___U13081 ( .A1(register__n12288), .A2(register__n1931), .B1(register__n9531), .B2(register__n1929), 
        .Y(register__n12870) );
  OA22x2_ASAP7_75t_R register___U13082 ( .A1(register__n3305), .A2(register__n893), .B1(register__n10434), .B2(register__n896), 
        .Y(register__n13056) );
  INVx1_ASAP7_75t_R register___U13083 ( .A(register__n5085), .Y(register__n8663) );
  OA22x2_ASAP7_75t_R register___U13084 ( .A1(register__net63244), .A2(register__n1140), .B1(register__net91263), .B2(
        n1144), .Y(register__n13154) );
  OA22x2_ASAP7_75t_R register___U13085 ( .A1(register__n12170), .A2(register__n118), .B1(register__n9561), .B2(register__n1190), 
        .Y(register__n13101) );
  OA22x2_ASAP7_75t_R register___U13086 ( .A1(register__n12110), .A2(register__n460), .B1(register__n9433), .B2(register__n467), 
        .Y(register__n12937) );
  OA22x2_ASAP7_75t_R register___U13087 ( .A1(register__n12279), .A2(register__n3719), .B1(register__n9563), .B2(register__n11848), 
        .Y(register__n13370) );
  BUFx12f_ASAP7_75t_R register___U13088 ( .A(register__net103542), .Y(register__net91219) );
  OA22x2_ASAP7_75t_R register___U13089 ( .A1(register__n12088), .A2(register__n2824), .B1(register__n9569), .B2(register__n1944), 
        .Y(register__n12878) );
  INVx1_ASAP7_75t_R register___U13090 ( .A(register__n3932), .Y(register__n8669) );
  OA22x2_ASAP7_75t_R register___U13091 ( .A1(register__n12089), .A2(register__n1069), .B1(register__n10428), .B2(register__n81), 
        .Y(register__n12822) );
  INVx1_ASAP7_75t_R register___U13092 ( .A(register__n6512), .Y(register__n8670) );
  OA22x2_ASAP7_75t_R register___U13093 ( .A1(register__register__n12023), .A2(register__n120), .B1(register__n10343), .B2(register__n1211), 
        .Y(register__n13112) );
  OA22x2_ASAP7_75t_R register___U13094 ( .A1(register__net64920), .A2(register__n1568), .B1(register__n10341), .B2(
        n1206), .Y(register__n13111) );
  INVx1_ASAP7_75t_R register___U13095 ( .A(register__n5793), .Y(register__n8671) );
  OA22x2_ASAP7_75t_R register___U13096 ( .A1(register__net64934), .A2(register__n109), .B1(register__n9961), .B2(register__n5838), 
        .Y(register__n12856) );
  OA22x2_ASAP7_75t_R register___U13097 ( .A1(register__n12199), .A2(register__n461), .B1(register__n9423), .B2(register__n468), 
        .Y(register__n12933) );
  INVx1_ASAP7_75t_R register___U13098 ( .A(register__n4773), .Y(register__n8674) );
  OA22x2_ASAP7_75t_R register___U13099 ( .A1(register__n12197), .A2(register__n889), .B1(register__n9409), .B2(register__n900), 
        .Y(register__n13050) );
  INVx1_ASAP7_75t_R register___U13100 ( .A(register__n5081), .Y(register__n8675) );
  OA22x2_ASAP7_75t_R register___U13101 ( .A1(register__n12149), .A2(register__n109), .B1(register__n10094), .B2(register__n6720), 
        .Y(register__n12847) );
  OA22x2_ASAP7_75t_R register___U13102 ( .A1(register__net62996), .A2(register__n953), .B1(register__n10442), .B2(register__n960), 
        .Y(register__n13013) );
  OA22x2_ASAP7_75t_R register___U13103 ( .A1(register__n12455), .A2(register__n1137), .B1(register__n10385), .B2(register__n1150), 
        .Y(register__n13149) );
  OA22x2_ASAP7_75t_R register___U13104 ( .A1(register__n12462), .A2(register__n176), .B1(register__n9796), .B2(register__n214), 
        .Y(register__n12662) );
  OA22x2_ASAP7_75t_R register___U13105 ( .A1(register__n12432), .A2(register__n190), .B1(register__n9343), .B2(register__n217), 
        .Y(register__n12664) );
  INVx1_ASAP7_75t_R register___U13106 ( .A(register__n12664), .Y(register__n8678) );
  OA22x2_ASAP7_75t_R register___U13107 ( .A1(register__n12459), .A2(register__n2827), .B1(register__n9525), .B2(register__n1887), 
        .Y(register__n12860) );
  INVx1_ASAP7_75t_R register___U13108 ( .A(register__n4076), .Y(register__n8679) );
  OA22x2_ASAP7_75t_R register___U13109 ( .A1(register__net62830), .A2(register__n1415), .B1(register__net90229), .B2(
        n1418), .Y(register__n12981) );
  OA22x2_ASAP7_75t_R register___U13110 ( .A1(register__n3304), .A2(register__n118), .B1(register__n10375), .B2(register__n1201), 
        .Y(register__n13090) );
  INVx1_ASAP7_75t_R register___U13111 ( .A(register__n4070), .Y(register__n8680) );
  OA22x2_ASAP7_75t_R register___U13112 ( .A1(register__net109773), .A2(register__n3343), .B1(register__n10501), .B2(
        n11780), .Y(register__n12950) );
  OA22x2_ASAP7_75t_R register___U13113 ( .A1(register__n12428), .A2(register__n461), .B1(register__n10136), .B2(register__n473), 
        .Y(register__n12922) );
  INVx1_ASAP7_75t_R register___U13114 ( .A(register__n3956), .Y(register__n8682) );
  OA22x2_ASAP7_75t_R register___U13115 ( .A1(register__n12461), .A2(register__n337), .B1(register__n9792), .B2(register__n343), 
        .Y(register__n12718) );
  OA22x2_ASAP7_75t_R register___U13116 ( .A1(register__n12427), .A2(register__n101), .B1(register__n9301), .B2(register__n2010), 
        .Y(register__n12952) );
  OA22x2_ASAP7_75t_R register___U13117 ( .A1(register__n12424), .A2(register__n103), .B1(register__register__n10395), .B2(register__n1147), 
        .Y(register__n13151) );
  OA22x2_ASAP7_75t_R register___U13118 ( .A1(register__net62826), .A2(register__n1120), .B1(register__net90237), .B2(
        n3476), .Y(register__n13065) );
  OR3x1_ASAP7_75t_R register___U13119 ( .A(register__n5451), .B(register__n8692), .C(register__n8690), .Y(register__n11221) );
  OA22x2_ASAP7_75t_R register___U13120 ( .A1(register__net131654), .A2(register__n7341), .B1(register__net130175), .B2(
        n10596), .Y(register__n11224) );
  INVx1_ASAP7_75t_R register___U13121 ( .A(register__n5449), .Y(register__n8690) );
  OA222x2_ASAP7_75t_R register___U13122 ( .A1(register__n1987), .A2(register__n10599), .B1(register__n1995), .B2(register__n10600), .C1(register__n1800), .C2(register__n6762), .Y(register__n11222) );
  OA22x2_ASAP7_75t_R register___U13123 ( .A1(register__n714), .A2(register__n7092), .B1(register__n10598), .B2(register__n407), 
        .Y(register__n11223) );
  INVx1_ASAP7_75t_R register___U13124 ( .A(register__n5452), .Y(register__n8692) );
  OR3x1_ASAP7_75t_R register___U13125 ( .A(register__n4755), .B(register__n8695), .C(register__n8694), .Y(register__n10591) );
  OA22x2_ASAP7_75t_R register___U13126 ( .A1(register__n420), .A2(register__register__n8003), .B1(register__n800), .B2(register__n6766), 
        .Y(register__n10594) );
  INVx1_ASAP7_75t_R register___U13127 ( .A(register__n4749), .Y(register__n8694) );
  OA22x2_ASAP7_75t_R register___U13128 ( .A1(register__net107674), .A2(register__n7339), .B1(register__n1691), .B2(
        n7688), .Y(register__n10593) );
  INVx1_ASAP7_75t_R register___U13129 ( .A(register__n4751), .Y(register__n8695) );
  OA222x2_ASAP7_75t_R register___U13130 ( .A1(register__n2002), .A2(register__n5730), .B1(register__n817), .B2(register__n6210), 
        .C1(register__net112580), .C2(register__n11227), .Y(register__n10592) );
  OR3x1_ASAP7_75t_R register___U13131 ( .A(register__n486), .B(register__n8699), .C(register__n8698), .Y(register__n10909) );
  OA22x2_ASAP7_75t_R register___U13132 ( .A1(register__n420), .A2(register__n6485), .B1(register__n800), .B2(register__n6230), 
        .Y(register__n10912) );
  INVx1_ASAP7_75t_R register___U13133 ( .A(register__n5134), .Y(register__n8698) );
  OA22x2_ASAP7_75t_R register___U13134 ( .A1(register__net107674), .A2(register__n11525), .B1(register__n1691), .B2(
        n7867), .Y(register__n10911) );
  INVx1_ASAP7_75t_R register___U13135 ( .A(register__n5136), .Y(register__n8699) );
  OR3x1_ASAP7_75t_R register___U13136 ( .A(register__n4951), .B(register__n8701), .C(register__n8700), .Y(register__n11056) );
  OA22x2_ASAP7_75t_R register___U13137 ( .A1(register__n420), .A2(register__n7106), .B1(register__n800), .B2(register__n11060), 
        .Y(register__n11058) );
  OA22x2_ASAP7_75t_R register___U13138 ( .A1(register__n66), .A2(register__n7696), .B1(register__n1691), .B2(register__n8007), 
        .Y(register__n11057) );
  INVx1_ASAP7_75t_R register___U13139 ( .A(register__n4949), .Y(register__n8701) );
  OR3x1_ASAP7_75t_R register___U13140 ( .A(register__n5819), .B(register__n8704), .C(register__n8703), .Y(register__n11387) );
  OA22x2_ASAP7_75t_R register___U13141 ( .A1(register__n1965), .A2(register__n11391), .B1(register__net130175), .B2(
        n7097), .Y(register__n11390) );
  INVx1_ASAP7_75t_R register___U13142 ( .A(register__n5813), .Y(register__n8703) );
  OA22x2_ASAP7_75t_R register___U13143 ( .A1(register__n712), .A2(register__n7344), .B1(register__n353), .B2(register__n8004), 
        .Y(register__n11389) );
  INVx1_ASAP7_75t_R register___U13144 ( .A(register__n5815), .Y(register__n8704) );
  INVx1_ASAP7_75t_R register___U13145 ( .A(register__n5817), .Y(register__n8705) );
  OA22x2_ASAP7_75t_R register___U13146 ( .A1(register__n2013), .A2(register__n7691), .B1(register__net130175), .B2(
        n6484), .Y(register__n11178) );
  INVx1_ASAP7_75t_R register___U13147 ( .A(register__n5806), .Y(register__n8744) );
  OA222x2_ASAP7_75t_R register___U13148 ( .A1(register__net127626), .A2(register__n10556), .B1(register__n1995), .B2(
        n6983), .C1(register__n1800), .C2(register__n6209), .Y(register__n11176) );
  OA22x2_ASAP7_75t_R register___U13149 ( .A1(register__n713), .A2(register__n5956), .B1(register__n353), .B2(register__n7244), 
        .Y(register__n11177) );
  INVx1_ASAP7_75t_R register___U13150 ( .A(register__n5811), .Y(register__n8746) );
  OR3x1_ASAP7_75t_R register___U13151 ( .A(register__n8750), .B(register__n8748), .C(register__n8749), .Y(register__n11122) );
  OA22x2_ASAP7_75t_R register___U13152 ( .A1(register__net107674), .A2(register__n7693), .B1(register__n1691), .B2(
        n11129), .Y(register__n11124) );
  INVx1_ASAP7_75t_R register___U13153 ( .A(register__n5153), .Y(register__n8748) );
  OA22x2_ASAP7_75t_R register___U13154 ( .A1(register__n420), .A2(register__n11126), .B1(register__n800), .B2(register__n11127), 
        .Y(register__n11125) );
  INVx1_ASAP7_75t_R register___U13155 ( .A(register__n5155), .Y(register__n8749) );
  OA222x2_ASAP7_75t_R register___U13156 ( .A1(register__n2002), .A2(register__n11130), .B1(register__n1997), .B2(
        C6423_net61304), .C1(register__net112580), .C2(register__n7576), .Y(register__n11123) );
  INVx1_ASAP7_75t_R register___U13157 ( .A(register__n11123), .Y(register__n8750) );
  OA22x2_ASAP7_75t_R register___U13158 ( .A1(register__n2013), .A2(register__n8006), .B1(register__net130175), .B2(
        n6231), .Y(register__n11453) );
  OA22x2_ASAP7_75t_R register___U13159 ( .A1(register__n711), .A2(register__n6780), .B1(register__net149934), .B2(register__n7242), .Y(register__n11452) );
  OA222x2_ASAP7_75t_R register___U13160 ( .A1(register__n1987), .A2(register__n6477), .B1(register__n1995), .B2(register__n11458), 
        .C1(register__n1800), .C2(register__n7575), .Y(register__n11451) );
  BUFx6f_ASAP7_75t_R register___U13161 ( .A(register__n8754), .Y(register__n8753) );
  BUFx4f_ASAP7_75t_R register___U13162 ( .A(register__n7497), .Y(register__n8754) );
  BUFx4f_ASAP7_75t_R register___U13163 ( .A(register__net109898), .Y(register__net96915) );
  BUFx6f_ASAP7_75t_R register___U13164 ( .A(register__n8756), .Y(register__n8755) );
  BUFx4f_ASAP7_75t_R register___U13165 ( .A(register__n5359), .Y(register__n8756) );
  BUFx6f_ASAP7_75t_R register___U13166 ( .A(register__n8758), .Y(register__n8757) );
  BUFx4f_ASAP7_75t_R register___U13167 ( .A(register__n6550), .Y(register__n8758) );
  BUFx4f_ASAP7_75t_R register___U13168 ( .A(register__net108071), .Y(register__net96903) );
  BUFx6f_ASAP7_75t_R register___U13169 ( .A(register__n8760), .Y(register__n8759) );
  BUFx4f_ASAP7_75t_R register___U13170 ( .A(register__n6088), .Y(register__n8760) );
  BUFx4f_ASAP7_75t_R register___U13171 ( .A(register__net108067), .Y(register__net96895) );
  BUFx6f_ASAP7_75t_R register___U13172 ( .A(register__n8762), .Y(register__n8761) );
  BUFx4f_ASAP7_75t_R register___U13173 ( .A(register__n6090), .Y(register__n8762) );
  BUFx6f_ASAP7_75t_R register___U13174 ( .A(register__n8764), .Y(register__n8763) );
  BUFx4f_ASAP7_75t_R register___U13175 ( .A(register__n7739), .Y(register__n8764) );
  BUFx6f_ASAP7_75t_R register___U13176 ( .A(register__n8766), .Y(register__n8765) );
  BUFx4f_ASAP7_75t_R register___U13177 ( .A(register__n6860), .Y(register__n8766) );
  BUFx6f_ASAP7_75t_R register___U13178 ( .A(register__n8768), .Y(register__n8767) );
  BUFx4f_ASAP7_75t_R register___U13179 ( .A(register__n7753), .Y(register__n8768) );
  BUFx6f_ASAP7_75t_R register___U13180 ( .A(register__n8770), .Y(register__n8769) );
  BUFx4f_ASAP7_75t_R register___U13181 ( .A(register__n6354), .Y(register__n8770) );
  BUFx6f_ASAP7_75t_R register___U13182 ( .A(register__n8772), .Y(register__n8771) );
  BUFx4f_ASAP7_75t_R register___U13183 ( .A(register__n3747), .Y(register__n8772) );
  BUFx6f_ASAP7_75t_R register___U13184 ( .A(register__n8774), .Y(register__n8773) );
  BUFx4f_ASAP7_75t_R register___U13185 ( .A(register__n6890), .Y(register__n8774) );
  BUFx4f_ASAP7_75t_R register___U13186 ( .A(register__net126192), .Y(register__net96863) );
  BUFx6f_ASAP7_75t_R register___U13187 ( .A(register__n8776), .Y(register__n8775) );
  BUFx4f_ASAP7_75t_R register___U13188 ( .A(register__n5887), .Y(register__n8776) );
  BUFx6f_ASAP7_75t_R register___U13189 ( .A(register__n8778), .Y(register__n8777) );
  BUFx4f_ASAP7_75t_R register___U13190 ( .A(register__n3749), .Y(register__n8778) );
  BUFx4f_ASAP7_75t_R register___U13191 ( .A(register__n8187), .Y(register__n8780) );
  BUFx6f_ASAP7_75t_R register___U13192 ( .A(register__n8782), .Y(register__n8781) );
  BUFx4f_ASAP7_75t_R register___U13193 ( .A(register__n6124), .Y(register__n8782) );
  BUFx4f_ASAP7_75t_R register___U13194 ( .A(register__net107852), .Y(register__net96843) );
  BUFx4f_ASAP7_75t_R register___U13195 ( .A(register__n5202), .Y(register__n8784) );
  BUFx6f_ASAP7_75t_R register___U13196 ( .A(register__n8786), .Y(register__n8785) );
  BUFx4f_ASAP7_75t_R register___U13197 ( .A(register__n6565), .Y(register__n8786) );
  BUFx6f_ASAP7_75t_R register___U13198 ( .A(register__n8788), .Y(register__n8787) );
  BUFx4f_ASAP7_75t_R register___U13199 ( .A(register__n6569), .Y(register__n8788) );
  BUFx6f_ASAP7_75t_R register___U13200 ( .A(register__n8790), .Y(register__n8789) );
  BUFx4f_ASAP7_75t_R register___U13201 ( .A(register__n3800), .Y(register__n8790) );
  BUFx6f_ASAP7_75t_R register___U13202 ( .A(register__n8792), .Y(register__n8791) );
  BUFx4f_ASAP7_75t_R register___U13203 ( .A(register__n7464), .Y(register__n8792) );
  BUFx4f_ASAP7_75t_R register___U13204 ( .A(register__net103552), .Y(register__net96819) );
  BUFx6f_ASAP7_75t_R register___U13205 ( .A(register__n8794), .Y(register__n8793) );
  BUFx4f_ASAP7_75t_R register___U13206 ( .A(register__n7223), .Y(register__n8794) );
  BUFx6f_ASAP7_75t_R register___U13207 ( .A(register__n8796), .Y(register__n8795) );
  BUFx4f_ASAP7_75t_R register___U13208 ( .A(register__n7408), .Y(register__n8796) );
  BUFx6f_ASAP7_75t_R register___U13209 ( .A(register__n8798), .Y(register__n8797) );
  BUFx4f_ASAP7_75t_R register___U13210 ( .A(register__n6101), .Y(register__n8798) );
  BUFx4f_ASAP7_75t_R register___U13211 ( .A(register__net110024), .Y(register__net96767) );
  BUFx6f_ASAP7_75t_R register___U13212 ( .A(register__n8800), .Y(register__n8799) );
  BUFx4f_ASAP7_75t_R register___U13213 ( .A(register__n7161), .Y(register__n8800) );
  BUFx6f_ASAP7_75t_R register___U13214 ( .A(register__n8802), .Y(register__n8801) );
  BUFx4f_ASAP7_75t_R register___U13215 ( .A(register__n8066), .Y(register__n8802) );
  BUFx4f_ASAP7_75t_R register___U13216 ( .A(register__n7854), .Y(register__n8804) );
  BUFx6f_ASAP7_75t_R register___U13217 ( .A(register__n8806), .Y(register__n8805) );
  BUFx4f_ASAP7_75t_R register___U13218 ( .A(register__n5847), .Y(register__n8806) );
  BUFx6f_ASAP7_75t_R register___U13219 ( .A(register__n8808), .Y(register__n8807) );
  BUFx4f_ASAP7_75t_R register___U13220 ( .A(register__n6334), .Y(register__n8808) );
  BUFx6f_ASAP7_75t_R register___U13221 ( .A(register__n8810), .Y(register__n8809) );
  BUFx4f_ASAP7_75t_R register___U13222 ( .A(register__n6103), .Y(register__n8810) );
  BUFx6f_ASAP7_75t_R register___U13223 ( .A(register__n8812), .Y(register__n8811) );
  BUFx4f_ASAP7_75t_R register___U13224 ( .A(register__n7187), .Y(register__n8812) );
  BUFx6f_ASAP7_75t_R register___U13225 ( .A(register__n8814), .Y(register__n8813) );
  BUFx4f_ASAP7_75t_R register___U13226 ( .A(register__n3697), .Y(register__n8814) );
  BUFx6f_ASAP7_75t_R register___U13227 ( .A(register__n8816), .Y(register__n8815) );
  BUFx4f_ASAP7_75t_R register___U13228 ( .A(register__n7567), .Y(register__n8816) );
  BUFx6f_ASAP7_75t_R register___U13229 ( .A(register__n8818), .Y(register__n8817) );
  BUFx4f_ASAP7_75t_R register___U13230 ( .A(register__n3794), .Y(register__n8818) );
  BUFx6f_ASAP7_75t_R register___U13231 ( .A(register__n8822), .Y(register__n8821) );
  BUFx4f_ASAP7_75t_R register___U13232 ( .A(register__n6386), .Y(register__n8822) );
  BUFx6f_ASAP7_75t_R register___U13233 ( .A(register__n8824), .Y(register__n8823) );
  BUFx4f_ASAP7_75t_R register___U13234 ( .A(register__n7218), .Y(register__n8824) );
  BUFx6f_ASAP7_75t_R register___U13235 ( .A(register__n8826), .Y(register__n8825) );
  BUFx4f_ASAP7_75t_R register___U13236 ( .A(register__n7443), .Y(register__n8826) );
  BUFx6f_ASAP7_75t_R register___U13237 ( .A(register__n8828), .Y(register__n8827) );
  BUFx4f_ASAP7_75t_R register___U13238 ( .A(register__n7743), .Y(register__n8828) );
  BUFx6f_ASAP7_75t_R register___U13239 ( .A(register__net96611), .Y(register__net96610) );
  BUFx4f_ASAP7_75t_R register___U13240 ( .A(register__net103708), .Y(register__net96611) );
  BUFx6f_ASAP7_75t_R register___U13241 ( .A(register__n8830), .Y(register__n8829) );
  BUFx4f_ASAP7_75t_R register___U13242 ( .A(register__n7813), .Y(register__n8830) );
  BUFx6f_ASAP7_75t_R register___U13243 ( .A(register__n8832), .Y(register__n8831) );
  BUFx4f_ASAP7_75t_R register___U13244 ( .A(register__n7824), .Y(register__n8832) );
  BUFx6f_ASAP7_75t_R register___U13245 ( .A(register__n8834), .Y(register__n8833) );
  BUFx4f_ASAP7_75t_R register___U13246 ( .A(register__n7835), .Y(register__n8834) );
  BUFx2_ASAP7_75t_R register___U13247 ( .A(register__n10639), .Y(register__n8837) );
  BUFx2_ASAP7_75t_R register___U13248 ( .A(Reg_data[116]), .Y(register__n8838) );
  BUFx12f_ASAP7_75t_R register___U13249 ( .A(register__n8840), .Y(register__n8839) );
  BUFx12f_ASAP7_75t_R register___U13250 ( .A(register__n10037), .Y(register__n8840) );
  BUFx12f_ASAP7_75t_R register___U13251 ( .A(register__n8839), .Y(register__n10036) );
  BUFx2_ASAP7_75t_R register___U13252 ( .A(Reg_data[49]), .Y(register__n8841) );
  BUFx12f_ASAP7_75t_R register___U13253 ( .A(register__n10121), .Y(register__n8842) );
  BUFx12f_ASAP7_75t_R register___U13254 ( .A(register__n8842), .Y(register__n10120) );
  BUFx4f_ASAP7_75t_R register___U13255 ( .A(register__n6811), .Y(register__n10121) );
  BUFx2_ASAP7_75t_R register___U13256 ( .A(Reg_data[110]), .Y(register__n8843) );
  BUFx12f_ASAP7_75t_R register___U13257 ( .A(register__n10141), .Y(register__n8844) );
  BUFx12f_ASAP7_75t_R register___U13258 ( .A(register__n8844), .Y(register__n10140) );
  BUFx2_ASAP7_75t_R register___U13259 ( .A(Reg_data[125]), .Y(register__net95809) );
  BUFx4f_ASAP7_75t_R register___U13260 ( .A(register__net98937), .Y(register__net89445) );
  BUFx3_ASAP7_75t_R register___U13261 ( .A(register__net95679), .Y(register__net95678) );
  BUFx2_ASAP7_75t_R register___U13262 ( .A(Reg_data[857]), .Y(register__net95679) );
  BUFx3_ASAP7_75t_R register___U13263 ( .A(register__n8846), .Y(register__n8845) );
  BUFx2_ASAP7_75t_R register___U13264 ( .A(Reg_data[848]), .Y(register__n8846) );
  BUFx3_ASAP7_75t_R register___U13265 ( .A(register__n8848), .Y(register__n8847) );
  BUFx2_ASAP7_75t_R register___U13266 ( .A(Reg_data[840]), .Y(register__n8848) );
  BUFx3_ASAP7_75t_R register___U13267 ( .A(register__n8850), .Y(register__n8849) );
  BUFx2_ASAP7_75t_R register___U13268 ( .A(Reg_data[835]), .Y(register__n8850) );
  BUFx3_ASAP7_75t_R register___U13269 ( .A(register__n8852), .Y(register__n8851) );
  BUFx2_ASAP7_75t_R register___U13270 ( .A(Reg_data[788]), .Y(register__n8852) );
  BUFx3_ASAP7_75t_R register___U13271 ( .A(register__n8854), .Y(register__n8853) );
  BUFx2_ASAP7_75t_R register___U13272 ( .A(Reg_data[776]), .Y(register__n8854) );
  BUFx3_ASAP7_75t_R register___U13273 ( .A(register__n8856), .Y(register__n8855) );
  BUFx2_ASAP7_75t_R register___U13274 ( .A(Reg_data[771]), .Y(register__n8856) );
  BUFx3_ASAP7_75t_R register___U13275 ( .A(register__n8858), .Y(register__n8857) );
  BUFx2_ASAP7_75t_R register___U13276 ( .A(Reg_data[769]), .Y(register__n8858) );
  BUFx3_ASAP7_75t_R register___U13277 ( .A(register__net95647), .Y(register__net95646) );
  BUFx2_ASAP7_75t_R register___U13278 ( .A(Reg_data[677]), .Y(register__net95647) );
  BUFx3_ASAP7_75t_R register___U13279 ( .A(register__n8860), .Y(register__n8859) );
  BUFx2_ASAP7_75t_R register___U13280 ( .A(Reg_data[675]), .Y(register__n8860) );
  BUFx3_ASAP7_75t_R register___U13281 ( .A(register__n8862), .Y(register__n8861) );
  BUFx2_ASAP7_75t_R register___U13282 ( .A(Reg_data[673]), .Y(register__n8862) );
  BUFx3_ASAP7_75t_R register___U13283 ( .A(register__n8864), .Y(register__n8863) );
  BUFx2_ASAP7_75t_R register___U13284 ( .A(Reg_data[596]), .Y(register__n8864) );
  BUFx3_ASAP7_75t_R register___U13285 ( .A(register__n8866), .Y(register__n8865) );
  BUFx2_ASAP7_75t_R register___U13286 ( .A(Reg_data[592]), .Y(register__n8866) );
  BUFx3_ASAP7_75t_R register___U13287 ( .A(register__n8868), .Y(register__n8867) );
  BUFx2_ASAP7_75t_R register___U13288 ( .A(Reg_data[579]), .Y(register__n8868) );
  BUFx3_ASAP7_75t_R register___U13289 ( .A(register__n8870), .Y(register__n8869) );
  BUFx2_ASAP7_75t_R register___U13290 ( .A(Reg_data[448]), .Y(register__n8870) );
  BUFx3_ASAP7_75t_R register___U13291 ( .A(register__net95619), .Y(register__net95618) );
  BUFx2_ASAP7_75t_R register___U13292 ( .A(Reg_data[441]), .Y(register__net95619) );
  BUFx3_ASAP7_75t_R register___U13293 ( .A(register__n8872), .Y(register__n8871) );
  BUFx2_ASAP7_75t_R register___U13294 ( .A(Reg_data[438]), .Y(register__n8872) );
  BUFx3_ASAP7_75t_R register___U13295 ( .A(register__n8874), .Y(register__n8873) );
  BUFx2_ASAP7_75t_R register___U13296 ( .A(Reg_data[385]), .Y(register__n8874) );
  BUFx3_ASAP7_75t_R register___U13297 ( .A(register__n8876), .Y(register__n8875) );
  BUFx2_ASAP7_75t_R register___U13298 ( .A(Reg_data[373]), .Y(register__n8876) );
  BUFx3_ASAP7_75t_R register___U13299 ( .A(register__n8878), .Y(register__n8877) );
  BUFx2_ASAP7_75t_R register___U13300 ( .A(Reg_data[372]), .Y(register__n8878) );
  BUFx3_ASAP7_75t_R register___U13301 ( .A(register__n8880), .Y(register__n8879) );
  BUFx2_ASAP7_75t_R register___U13302 ( .A(Reg_data[370]), .Y(register__n8880) );
  BUFx3_ASAP7_75t_R register___U13303 ( .A(register__net95595), .Y(register__net95594) );
  BUFx2_ASAP7_75t_R register___U13304 ( .A(Reg_data[357]), .Y(register__net95595) );
  BUFx3_ASAP7_75t_R register___U13305 ( .A(register__n8882), .Y(register__n8881) );
  BUFx2_ASAP7_75t_R register___U13306 ( .A(Reg_data[340]), .Y(register__n8882) );
  BUFx3_ASAP7_75t_R register___U13307 ( .A(register__n8884), .Y(register__n8883) );
  BUFx2_ASAP7_75t_R register___U13308 ( .A(Reg_data[324]), .Y(register__n8884) );
  BUFx3_ASAP7_75t_R register___U13309 ( .A(register__n8886), .Y(register__n8885) );
  BUFx2_ASAP7_75t_R register___U13310 ( .A(Reg_data[323]), .Y(register__n8886) );
  BUFx3_ASAP7_75t_R register___U13311 ( .A(register__n8888), .Y(register__n8887) );
  BUFx2_ASAP7_75t_R register___U13312 ( .A(Reg_data[259]), .Y(register__n8888) );
  BUFx3_ASAP7_75t_R register___U13313 ( .A(register__net95572), .Y(register__net95571) );
  BUFx2_ASAP7_75t_R register___U13314 ( .A(Reg_data[121]), .Y(register__net95572) );
  BUFx12f_ASAP7_75t_R register___U13315 ( .A(register__net101570), .Y(register__net89845) );
  BUFx3_ASAP7_75t_R register___U13316 ( .A(register__n8890), .Y(register__n8889) );
  BUFx2_ASAP7_75t_R register___U13317 ( .A(Reg_data[117]), .Y(register__n8890) );
  BUFx12f_ASAP7_75t_R register___U13318 ( .A(register__n10035), .Y(register__n8891) );
  BUFx12f_ASAP7_75t_R register___U13319 ( .A(register__n8891), .Y(register__n10034) );
  BUFx3_ASAP7_75t_R register___U13320 ( .A(register__net95558), .Y(register__net95557) );
  BUFx2_ASAP7_75t_R register___U13321 ( .A(Reg_data[101]), .Y(register__net95558) );
  BUFx12f_ASAP7_75t_R register___U13322 ( .A(register__net89814), .Y(register__net89813) );
  BUFx3_ASAP7_75t_R register___U13323 ( .A(register__n8893), .Y(register__n8892) );
  BUFx2_ASAP7_75t_R register___U13324 ( .A(Reg_data[100]), .Y(register__n8893) );
  BUFx12f_ASAP7_75t_R register___U13325 ( .A(register__n10045), .Y(register__n8894) );
  BUFx12f_ASAP7_75t_R register___U13326 ( .A(register__n8894), .Y(register__n10044) );
  BUFx3_ASAP7_75t_R register___U13327 ( .A(register__n8896), .Y(register__n8895) );
  BUFx2_ASAP7_75t_R register___U13328 ( .A(Reg_data[97]), .Y(register__n8896) );
  BUFx12f_ASAP7_75t_R register___U13329 ( .A(register__n8898), .Y(register__n8897) );
  BUFx12f_ASAP7_75t_R register___U13330 ( .A(register__n10455), .Y(register__n8898) );
  BUFx12f_ASAP7_75t_R register___U13331 ( .A(register__n8897), .Y(register__n10454) );
  BUFx3_ASAP7_75t_R register___U13332 ( .A(register__n8900), .Y(register__n8899) );
  BUFx2_ASAP7_75t_R register___U13333 ( .A(Reg_data[96]), .Y(register__n8900) );
  BUFx12f_ASAP7_75t_R register___U13334 ( .A(register__n10051), .Y(register__n8901) );
  BUFx12f_ASAP7_75t_R register___U13335 ( .A(register__n8901), .Y(register__n10050) );
  BUFx3_ASAP7_75t_R register___U13336 ( .A(register__n8903), .Y(register__n8902) );
  BUFx2_ASAP7_75t_R register___U13337 ( .A(Reg_data[84]), .Y(register__n8903) );
  BUFx3_ASAP7_75t_R register___U13338 ( .A(register__n8905), .Y(register__n8904) );
  BUFx2_ASAP7_75t_R register___U13339 ( .A(Reg_data[80]), .Y(register__n8905) );
  BUFx3_ASAP7_75t_R register___U13340 ( .A(register__n8907), .Y(register__n8906) );
  BUFx2_ASAP7_75t_R register___U13341 ( .A(Reg_data[67]), .Y(register__n8907) );
  BUFx3_ASAP7_75t_R register___U13342 ( .A(register__n8909), .Y(register__n8908) );
  BUFx2_ASAP7_75t_R register___U13343 ( .A(Reg_data[866]), .Y(register__n8909) );
  BUFx2_ASAP7_75t_R register___U13344 ( .A(register__n9698), .Y(register__n8910) );
  BUFx2_ASAP7_75t_R register___U13345 ( .A(register__n9698), .Y(register__n8911) );
  BUFx4f_ASAP7_75t_R register___U13346 ( .A(register__n9698), .Y(register__n8912) );
  BUFx3_ASAP7_75t_R register___U13347 ( .A(register__n8914), .Y(register__n8913) );
  BUFx2_ASAP7_75t_R register___U13348 ( .A(Reg_data[864]), .Y(register__n8914) );
  BUFx12f_ASAP7_75t_R register___U13349 ( .A(register__n9701), .Y(register__n8915) );
  BUFx12f_ASAP7_75t_R register___U13350 ( .A(register__n8915), .Y(register__n9700) );
  BUFx3_ASAP7_75t_R register___U13351 ( .A(register__net95499), .Y(register__net95498) );
  BUFx2_ASAP7_75t_R register___U13352 ( .A(Reg_data[889]), .Y(register__net95499) );
  BUFx12f_ASAP7_75t_R register___U13353 ( .A(register__net90762), .Y(register__net90761) );
  BUFx3_ASAP7_75t_R register___U13354 ( .A(register__n8917), .Y(register__n8916) );
  BUFx2_ASAP7_75t_R register___U13355 ( .A(Reg_data[886]), .Y(register__n8917) );
  BUFx3_ASAP7_75t_R register___U13356 ( .A(register__n8919), .Y(register__n8918) );
  BUFx2_ASAP7_75t_R register___U13357 ( .A(Reg_data[885]), .Y(register__n8919) );
  BUFx12f_ASAP7_75t_R register___U13358 ( .A(register__n9705), .Y(register__n8920) );
  BUFx12f_ASAP7_75t_R register___U13359 ( .A(register__n8920), .Y(register__n9704) );
  BUFx3_ASAP7_75t_R register___U13360 ( .A(register__n8922), .Y(register__n8921) );
  BUFx2_ASAP7_75t_R register___U13361 ( .A(Reg_data[865]), .Y(register__n8922) );
  BUFx12f_ASAP7_75t_R register___U13362 ( .A(register__n10500), .Y(register__n8923) );
  BUFx12f_ASAP7_75t_R register___U13363 ( .A(register__n8923), .Y(register__n10499) );
  BUFx3_ASAP7_75t_R register___U13364 ( .A(register__n8925), .Y(register__n8924) );
  BUFx2_ASAP7_75t_R register___U13365 ( .A(Reg_data[884]), .Y(register__n8925) );
  BUFx12f_ASAP7_75t_R register___U13366 ( .A(register__n8368), .Y(register__n8926) );
  BUFx12f_ASAP7_75t_R register___U13367 ( .A(register__n8926), .Y(register__n9706) );
  BUFx3_ASAP7_75t_R register___U13368 ( .A(register__n8928), .Y(register__n8927) );
  BUFx2_ASAP7_75t_R register___U13369 ( .A(Reg_data[882]), .Y(register__n8928) );
  BUFx2_ASAP7_75t_R register___U13370 ( .A(register__n9708), .Y(register__n8929) );
  BUFx2_ASAP7_75t_R register___U13371 ( .A(register__n9708), .Y(register__n8930) );
  BUFx4f_ASAP7_75t_R register___U13372 ( .A(register__n9708), .Y(register__n8931) );
  BUFx3_ASAP7_75t_R register___U13373 ( .A(register__n8933), .Y(register__n8932) );
  BUFx2_ASAP7_75t_R register___U13374 ( .A(Reg_data[880]), .Y(register__n8933) );
  BUFx3_ASAP7_75t_R register___U13375 ( .A(register__net95450), .Y(register__net95449) );
  BUFx2_ASAP7_75t_R register___U13376 ( .A(Reg_data[870]), .Y(register__net95450) );
  BUFx2_ASAP7_75t_R register___U13377 ( .A(register__net90733), .Y(register__net95451) );
  BUFx4f_ASAP7_75t_R register___U13378 ( .A(register__net90733), .Y(register__net95453) );
  BUFx3_ASAP7_75t_R register___U13379 ( .A(register__net95443), .Y(register__net95442) );
  BUFx2_ASAP7_75t_R register___U13380 ( .A(Reg_data[869]), .Y(register__net95443) );
  BUFx12f_ASAP7_75t_R register___U13381 ( .A(register__net90730), .Y(register__net90729) );
  BUFx3_ASAP7_75t_R register___U13382 ( .A(register__n8935), .Y(register__n8934) );
  BUFx2_ASAP7_75t_R register___U13383 ( .A(Reg_data[868]), .Y(register__n8935) );
  BUFx12f_ASAP7_75t_R register___U13384 ( .A(register__n9715), .Y(register__n8936) );
  BUFx12f_ASAP7_75t_R register___U13385 ( .A(register__n8936), .Y(register__n9714) );
  BUFx4f_ASAP7_75t_R register___U13386 ( .A(register__n8369), .Y(register__n8937) );
  BUFx2_ASAP7_75t_R register___U13387 ( .A(Reg_data[4]), .Y(register__n8938) );
  BUFx12f_ASAP7_75t_R register___U13388 ( .A(register__n8940), .Y(register__n8939) );
  BUFx12f_ASAP7_75t_R register___U13389 ( .A(register__n10356), .Y(register__n8940) );
  BUFx12f_ASAP7_75t_R register___U13390 ( .A(register__n8939), .Y(register__n10355) );
  BUFx6f_ASAP7_75t_R register___U13391 ( .A(register__n8937), .Y(register__n10356) );
  BUFx3_ASAP7_75t_R register___U13392 ( .A(register__n8942), .Y(register__n8941) );
  BUFx2_ASAP7_75t_R register___U13393 ( .A(Reg_data[3]), .Y(register__n8942) );
  BUFx3_ASAP7_75t_R register___U13394 ( .A(register__n8944), .Y(register__n8943) );
  BUFx2_ASAP7_75t_R register___U13395 ( .A(Reg_data[34]), .Y(register__n8944) );
  BUFx4f_ASAP7_75t_R register___U13396 ( .A(register__n10064), .Y(register__n8945) );
  BUFx2_ASAP7_75t_R register___U13397 ( .A(register__n10064), .Y(register__n8946) );
  BUFx2_ASAP7_75t_R register___U13398 ( .A(register__n10064), .Y(register__n8947) );
  BUFx3_ASAP7_75t_R register___U13399 ( .A(register__n8949), .Y(register__n8948) );
  BUFx2_ASAP7_75t_R register___U13400 ( .A(Reg_data[226]), .Y(register__n8949) );
  BUFx3_ASAP7_75t_R register___U13401 ( .A(register__n8951), .Y(register__n8950) );
  BUFx2_ASAP7_75t_R register___U13402 ( .A(Reg_data[54]), .Y(register__n8951) );
  BUFx12f_ASAP7_75t_R register___U13403 ( .A(register__n10073), .Y(register__n8952) );
  BUFx12f_ASAP7_75t_R register___U13404 ( .A(register__n8952), .Y(register__n10072) );
  BUFx3_ASAP7_75t_R register___U13405 ( .A(register__n8954), .Y(register__n8953) );
  BUFx2_ASAP7_75t_R register___U13406 ( .A(Reg_data[225]), .Y(register__n8954) );
  BUFx12f_ASAP7_75t_R register___U13407 ( .A(register__n10461), .Y(register__n8955) );
  BUFx12f_ASAP7_75t_R register___U13408 ( .A(register__n8955), .Y(register__n10460) );
  BUFx3_ASAP7_75t_R register___U13409 ( .A(register__n8957), .Y(register__n8956) );
  BUFx2_ASAP7_75t_R register___U13410 ( .A(Reg_data[52]), .Y(register__n8957) );
  BUFx12f_ASAP7_75t_R register___U13411 ( .A(register__n10079), .Y(register__n8958) );
  BUFx12f_ASAP7_75t_R register___U13412 ( .A(register__n8958), .Y(register__n10078) );
  BUFx3_ASAP7_75t_R register___U13413 ( .A(register__n8960), .Y(register__n8959) );
  BUFx2_ASAP7_75t_R register___U13414 ( .A(Reg_data[50]), .Y(register__n8960) );
  BUFx12f_ASAP7_75t_R register___U13415 ( .A(register__n10081), .Y(register__n8961) );
  BUFx12f_ASAP7_75t_R register___U13416 ( .A(register__n8961), .Y(register__n10080) );
  BUFx3_ASAP7_75t_R register___U13417 ( .A(register__net95373), .Y(register__net95372) );
  BUFx2_ASAP7_75t_R register___U13418 ( .A(Reg_data[37]), .Y(register__net95373) );
  BUFx12f_ASAP7_75t_R register___U13419 ( .A(register__net89714), .Y(register__net89713) );
  BUFx3_ASAP7_75t_R register___U13420 ( .A(register__net95366), .Y(register__net95365) );
  BUFx2_ASAP7_75t_R register___U13421 ( .A(Reg_data[229]), .Y(register__net95366) );
  BUFx2_ASAP7_75t_R register___U13422 ( .A(Reg_data[227]), .Y(register__n8963) );
  BUFx4f_ASAP7_75t_R register___U13423 ( .A(register__net101568), .Y(register__net95350) );
  BUFx2_ASAP7_75t_R register___U13424 ( .A(Reg_data[811]), .Y(register__net95351) );
  BUFx12f_ASAP7_75t_R register___U13425 ( .A(register__net90714), .Y(register__net90713) );
  BUFx6f_ASAP7_75t_R register___U13426 ( .A(register__net95350), .Y(register__net90714) );
  BUFx3_ASAP7_75t_R register___U13427 ( .A(register__net95341), .Y(register__net95340) );
  BUFx2_ASAP7_75t_R register___U13428 ( .A(Reg_data[907]), .Y(register__net95341) );
  BUFx3_ASAP7_75t_R register___U13429 ( .A(register__net88604), .Y(register__net95342) );
  BUFx4f_ASAP7_75t_R register___U13430 ( .A(register__net88604), .Y(register__net95344) );
  BUFx3_ASAP7_75t_R register___U13431 ( .A(register__n8965), .Y(register__n8964) );
  BUFx2_ASAP7_75t_R register___U13432 ( .A(Reg_data[781]), .Y(register__n8965) );
  BUFx4f_ASAP7_75t_R register___U13433 ( .A(register__n8016), .Y(register__n8966) );
  BUFx2_ASAP7_75t_R register___U13434 ( .A(Reg_data[103]), .Y(register__n8967) );
  BUFx12f_ASAP7_75t_R register___U13435 ( .A(register__n10097), .Y(register__n8968) );
  BUFx12f_ASAP7_75t_R register___U13436 ( .A(register__n8968), .Y(register__n10096) );
  BUFx6f_ASAP7_75t_R register___U13437 ( .A(register__n8966), .Y(register__n10097) );
  BUFx3_ASAP7_75t_R register___U13438 ( .A(register__net95322), .Y(register__net95321) );
  BUFx2_ASAP7_75t_R register___U13439 ( .A(Reg_data[619]), .Y(register__net95322) );
  BUFx12f_ASAP7_75t_R register___U13440 ( .A(register__net89662), .Y(register__net89661) );
  BUFx3_ASAP7_75t_R register___U13441 ( .A(register__n8970), .Y(register__n8969) );
  BUFx2_ASAP7_75t_R register___U13442 ( .A(Reg_data[269]), .Y(register__n8970) );
  BUFx3_ASAP7_75t_R register___U13443 ( .A(register__net95311), .Y(register__net95310) );
  BUFx2_ASAP7_75t_R register___U13444 ( .A(Reg_data[43]), .Y(register__net95311) );
  BUFx12f_ASAP7_75t_R register___U13445 ( .A(register__net89658), .Y(register__net89657) );
  BUFx3_ASAP7_75t_R register___U13446 ( .A(register__n8972), .Y(register__n8971) );
  BUFx2_ASAP7_75t_R register___U13447 ( .A(Reg_data[881]), .Y(register__n8972) );
  BUFx12f_ASAP7_75t_R register___U13448 ( .A(register__n9725), .Y(register__n8973) );
  BUFx12f_ASAP7_75t_R register___U13449 ( .A(register__n8973), .Y(register__n9724) );
  BUFx3_ASAP7_75t_R register___U13450 ( .A(register__n8975), .Y(register__n8974) );
  BUFx2_ASAP7_75t_R register___U13451 ( .A(Reg_data[589]), .Y(register__n8975) );
  BUFx3_ASAP7_75t_R register___U13452 ( .A(register__n8977), .Y(register__n8976) );
  BUFx2_ASAP7_75t_R register___U13453 ( .A(Reg_data[775]), .Y(register__n8977) );
  BUFx12f_ASAP7_75t_R register___U13454 ( .A(register__n8981), .Y(register__n8980) );
  BUFx12f_ASAP7_75t_R register___U13455 ( .A(register__n8980), .Y(register__n9513) );
  BUFx6f_ASAP7_75t_R register___U13456 ( .A(register__n8978), .Y(register__n9514) );
  BUFx3_ASAP7_75t_R register___U13457 ( .A(register__n8983), .Y(register__n8982) );
  BUFx2_ASAP7_75t_R register___U13458 ( .A(Reg_data[359]), .Y(register__n8983) );
  BUFx4f_ASAP7_75t_R register___U13459 ( .A(register__net101564), .Y(register__net95273) );
  BUFx2_ASAP7_75t_R register___U13460 ( .A(Reg_data[879]), .Y(register__net95274) );
  BUFx12f_ASAP7_75t_R register___U13461 ( .A(register__net90690), .Y(register__net90689) );
  BUFx6f_ASAP7_75t_R register___U13462 ( .A(register__net95273), .Y(register__net90690) );
  BUFx3_ASAP7_75t_R register___U13463 ( .A(register__n8985), .Y(register__n8984) );
  BUFx2_ASAP7_75t_R register___U13464 ( .A(Reg_data[607]), .Y(register__n8985) );
  BUFx4f_ASAP7_75t_R register___U13465 ( .A(register__n8371), .Y(register__n8986) );
  BUFx2_ASAP7_75t_R register___U13466 ( .A(Reg_data[109]), .Y(register__n8987) );
  BUFx12f_ASAP7_75t_R register___U13467 ( .A(register__n10109), .Y(register__n8988) );
  BUFx12f_ASAP7_75t_R register___U13468 ( .A(register__n8988), .Y(register__n10108) );
  BUFx6f_ASAP7_75t_R register___U13469 ( .A(register__n8986), .Y(register__n10109) );
  BUFx4f_ASAP7_75t_R register___U13470 ( .A(register__n8017), .Y(register__n8989) );
  BUFx2_ASAP7_75t_R register___U13471 ( .A(Reg_data[849]), .Y(register__n8990) );
  BUFx12f_ASAP7_75t_R register___U13472 ( .A(register__n8992), .Y(register__n8991) );
  BUFx12f_ASAP7_75t_R register___U13473 ( .A(register__n9518), .Y(register__n8992) );
  BUFx12f_ASAP7_75t_R register___U13474 ( .A(register__n8991), .Y(register__n9517) );
  BUFx6f_ASAP7_75t_R register___U13475 ( .A(register__n8989), .Y(register__n9518) );
  BUFx3_ASAP7_75t_R register___U13476 ( .A(register__net95242), .Y(register__net95241) );
  BUFx2_ASAP7_75t_R register___U13477 ( .A(Reg_data[875]), .Y(register__net95242) );
  BUFx4f_ASAP7_75t_R register___U13478 ( .A(register__net90677), .Y(register__net95245) );
  BUFx3_ASAP7_75t_R register___U13479 ( .A(register__net95235), .Y(register__net95234) );
  BUFx2_ASAP7_75t_R register___U13480 ( .A(Reg_data[363]), .Y(register__net95235) );
  BUFx12f_ASAP7_75t_R register___U13481 ( .A(register__net90670), .Y(register__net90669) );
  BUFx3_ASAP7_75t_R register___U13482 ( .A(register__net95228), .Y(register__net95227) );
  BUFx2_ASAP7_75t_R register___U13483 ( .A(Reg_data[683]), .Y(register__net95228) );
  BUFx12f_ASAP7_75t_R register___U13484 ( .A(register__net112724), .Y(register__net89597) );
  BUFx3_ASAP7_75t_R register___U13485 ( .A(register__net95221), .Y(register__net95220) );
  BUFx2_ASAP7_75t_R register___U13486 ( .A(Reg_data[235]), .Y(register__net95221) );
  BUFx12f_ASAP7_75t_R register___U13487 ( .A(register__net89582), .Y(register__net89581) );
  BUFx3_ASAP7_75t_R register___U13488 ( .A(register__n8994), .Y(register__n8993) );
  BUFx2_ASAP7_75t_R register___U13489 ( .A(Reg_data[327]), .Y(register__n8994) );
  BUFx4f_ASAP7_75t_R register___U13490 ( .A(register__n7374), .Y(register__n8995) );
  BUFx2_ASAP7_75t_R register___U13491 ( .A(Reg_data[890]), .Y(register__n8996) );
  BUFx12f_ASAP7_75t_R register___U13492 ( .A(register__n9733), .Y(register__n8997) );
  BUFx12f_ASAP7_75t_R register___U13493 ( .A(register__n8997), .Y(register__n9732) );
  BUFx6f_ASAP7_75t_R register___U13494 ( .A(register__n8995), .Y(register__n9733) );
  BUFx4f_ASAP7_75t_R register___U13495 ( .A(register__n8018), .Y(register__n8998) );
  BUFx12f_ASAP7_75t_R register___U13496 ( .A(register__n9001), .Y(register__n9000) );
  BUFx12f_ASAP7_75t_R register___U13497 ( .A(register__n9524), .Y(register__n9001) );
  BUFx12f_ASAP7_75t_R register___U13498 ( .A(register__n9000), .Y(register__n9523) );
  BUFx6f_ASAP7_75t_R register___U13499 ( .A(register__n8998), .Y(register__n9524) );
  BUFx3_ASAP7_75t_R register___U13500 ( .A(register__net95195), .Y(register__net95194) );
  BUFx2_ASAP7_75t_R register___U13501 ( .A(Reg_data[847]), .Y(register__net95195) );
  BUFx4f_ASAP7_75t_R register___U13502 ( .A(register__n8019), .Y(register__n9002) );
  BUFx2_ASAP7_75t_R register___U13503 ( .A(Reg_data[876]), .Y(register__n9003) );
  BUFx12f_ASAP7_75t_R register___U13504 ( .A(register__n9739), .Y(register__n9004) );
  BUFx12f_ASAP7_75t_R register___U13505 ( .A(register__n9004), .Y(register__n9738) );
  BUFx6f_ASAP7_75t_R register___U13506 ( .A(register__n9002), .Y(register__n9739) );
  BUFx3_ASAP7_75t_R register___U13507 ( .A(register__n9006), .Y(register__n9005) );
  BUFx2_ASAP7_75t_R register___U13508 ( .A(Reg_data[877]), .Y(register__n9006) );
  BUFx12f_ASAP7_75t_R register___U13509 ( .A(register__n9749), .Y(register__n9007) );
  BUFx12f_ASAP7_75t_R register___U13510 ( .A(register__n9007), .Y(register__n9748) );
  BUFx3_ASAP7_75t_R register___U13511 ( .A(register__n9009), .Y(register__n9008) );
  BUFx2_ASAP7_75t_R register___U13512 ( .A(Reg_data[333]), .Y(register__n9009) );
  BUFx3_ASAP7_75t_R register___U13513 ( .A(register__n9011), .Y(register__n9010) );
  BUFx2_ASAP7_75t_R register___U13514 ( .A(Reg_data[791]), .Y(register__n9011) );
  BUFx3_ASAP7_75t_R register___U13515 ( .A(register__n9013), .Y(register__n9012) );
  BUFx2_ASAP7_75t_R register___U13516 ( .A(Reg_data[602]), .Y(register__n9013) );
  BUFx4f_ASAP7_75t_R register___U13517 ( .A(register__n8020), .Y(register__n9014) );
  BUFx2_ASAP7_75t_R register___U13518 ( .A(Reg_data[119]), .Y(register__n9015) );
  BUFx12f_ASAP7_75t_R register___U13519 ( .A(register__n10129), .Y(register__n9016) );
  BUFx12f_ASAP7_75t_R register___U13520 ( .A(register__n9016), .Y(register__n10128) );
  BUFx6f_ASAP7_75t_R register___U13521 ( .A(register__n9014), .Y(register__n10129) );
  BUFx3_ASAP7_75t_R register___U13522 ( .A(register__n9018), .Y(register__n9017) );
  BUFx2_ASAP7_75t_R register___U13523 ( .A(Reg_data[671]), .Y(register__n9018) );
  BUFx3_ASAP7_75t_R register___U13524 ( .A(register__n9020), .Y(register__n9019) );
  BUFx2_ASAP7_75t_R register___U13525 ( .A(Reg_data[615]), .Y(register__n9020) );
  BUFx12f_ASAP7_75t_R register___U13526 ( .A(register__n10156), .Y(register__n9021) );
  BUFx12f_ASAP7_75t_R register___U13527 ( .A(register__n9021), .Y(register__n10155) );
  BUFx3_ASAP7_75t_R register___U13528 ( .A(register__n9023), .Y(register__n9022) );
  BUFx2_ASAP7_75t_R register___U13529 ( .A(Reg_data[17]), .Y(register__n9023) );
  BUFx3_ASAP7_75t_R register___U13530 ( .A(register__n9025), .Y(register__n9024) );
  BUFx2_ASAP7_75t_R register___U13531 ( .A(Reg_data[39]), .Y(register__n9025) );
  BUFx12f_ASAP7_75t_R register___U13532 ( .A(register__n7129), .Y(register__n9026) );
  BUFx12f_ASAP7_75t_R register___U13533 ( .A(register__n9026), .Y(register__n10160) );
  BUFx2_ASAP7_75t_R register___U13534 ( .A(Reg_data[231]), .Y(register__n9028) );
  BUFx3_ASAP7_75t_R register___U13535 ( .A(register__n9030), .Y(register__n9029) );
  BUFx2_ASAP7_75t_R register___U13536 ( .A(Reg_data[343]), .Y(register__n9030) );
  BUFx3_ASAP7_75t_R register___U13537 ( .A(register__n9032), .Y(register__n9031) );
  BUFx2_ASAP7_75t_R register___U13538 ( .A(Reg_data[858]), .Y(register__n9032) );
  BUFx3_ASAP7_75t_R register___U13539 ( .A(register__net95119), .Y(register__net95118) );
  BUFx2_ASAP7_75t_R register___U13540 ( .A(Reg_data[15]), .Y(register__net95119) );
  BUFx3_ASAP7_75t_R register___U13541 ( .A(register__net95115), .Y(register__net95114) );
  BUFx2_ASAP7_75t_R register___U13542 ( .A(Reg_data[285]), .Y(register__net95115) );
  BUFx3_ASAP7_75t_R register___U13543 ( .A(register__n9034), .Y(register__n9033) );
  BUFx2_ASAP7_75t_R register___U13544 ( .A(Reg_data[817]), .Y(register__n9034) );
  BUFx12f_ASAP7_75t_R register___U13545 ( .A(register__n9771), .Y(register__n9035) );
  BUFx12f_ASAP7_75t_R register___U13546 ( .A(register__n9035), .Y(register__n9770) );
  BUFx4f_ASAP7_75t_R register___U13547 ( .A(register__n8372), .Y(register__n9036) );
  BUFx2_ASAP7_75t_R register___U13548 ( .A(Reg_data[873]), .Y(register__n9037) );
  BUFx12f_ASAP7_75t_R register___U13549 ( .A(register__n9775), .Y(register__n9038) );
  BUFx12f_ASAP7_75t_R register___U13550 ( .A(register__n9038), .Y(register__n9774) );
  BUFx6f_ASAP7_75t_R register___U13551 ( .A(register__n9036), .Y(register__n9775) );
  BUFx3_ASAP7_75t_R register___U13552 ( .A(register__n9040), .Y(register__n9039) );
  BUFx2_ASAP7_75t_R register___U13553 ( .A(Reg_data[87]), .Y(register__n9040) );
  BUFx4f_ASAP7_75t_R register___U13554 ( .A(register__n5834), .Y(register__n9041) );
  BUFx2_ASAP7_75t_R register___U13555 ( .A(Reg_data[572]), .Y(register__n9042) );
  BUFx6f_ASAP7_75t_R register___U13556 ( .A(register__n9041), .Y(register__n10425) );
  BUFx3_ASAP7_75t_R register___U13557 ( .A(register__n9044), .Y(register__n9043) );
  BUFx2_ASAP7_75t_R register___U13558 ( .A(Reg_data[113]), .Y(register__n9044) );
  BUFx12f_ASAP7_75t_R register___U13559 ( .A(register__n10176), .Y(register__n9045) );
  BUFx12f_ASAP7_75t_R register___U13560 ( .A(register__n9045), .Y(register__n10175) );
  BUFx3_ASAP7_75t_R register___U13561 ( .A(register__net95071), .Y(register__net95070) );
  BUFx2_ASAP7_75t_R register___U13562 ( .A(Reg_data[239]), .Y(register__net95071) );
  BUFx2_ASAP7_75t_R register___U13563 ( .A(register__net91591), .Y(register__net95073) );
  BUFx3_ASAP7_75t_R register___U13564 ( .A(register__net95064), .Y(register__net95063) );
  BUFx2_ASAP7_75t_R register___U13565 ( .A(Reg_data[111]), .Y(register__net95064) );
  BUFx12f_ASAP7_75t_R register___U13566 ( .A(register__net89390), .Y(register__net89389) );
  BUFx3_ASAP7_75t_R register___U13567 ( .A(register__n9047), .Y(register__n9046) );
  BUFx2_ASAP7_75t_R register___U13568 ( .A(Reg_data[282]), .Y(register__n9047) );
  BUFx3_ASAP7_75t_R register___U13569 ( .A(register__n9049), .Y(register__n9048) );
  BUFx2_ASAP7_75t_R register___U13570 ( .A(Reg_data[871]), .Y(register__n9049) );
  BUFx12f_ASAP7_75t_R register___U13571 ( .A(register__n7707), .Y(register__n9050) );
  BUFx12f_ASAP7_75t_R register___U13572 ( .A(register__n9050), .Y(register__n9780) );
  BUFx3_ASAP7_75t_R register___U13573 ( .A(register__net95049), .Y(register__net95048) );
  BUFx2_ASAP7_75t_R register___U13574 ( .A(Reg_data[93]), .Y(register__net95049) );
  BUFx3_ASAP7_75t_R register___U13575 ( .A(register__n9052), .Y(register__n9051) );
  BUFx2_ASAP7_75t_R register___U13576 ( .A(Reg_data[894]), .Y(register__n9052) );
  BUFx3_ASAP7_75t_R register___U13577 ( .A(register__n9057), .Y(register__n9056) );
  BUFx2_ASAP7_75t_R register___U13578 ( .A(Reg_data[878]), .Y(register__n9057) );
  BUFx12f_ASAP7_75t_R register___U13579 ( .A(register__n7708), .Y(register__n9058) );
  BUFx12f_ASAP7_75t_R register___U13580 ( .A(register__n9058), .Y(register__n9802) );
  BUFx3_ASAP7_75t_R register___U13581 ( .A(register__n9060), .Y(register__n9059) );
  BUFx2_ASAP7_75t_R register___U13582 ( .A(Reg_data[734]), .Y(register__n9060) );
  BUFx4f_ASAP7_75t_R register___U13583 ( .A(register__n10219), .Y(register__n9061) );
  BUFx2_ASAP7_75t_R register___U13584 ( .A(register__n10219), .Y(register__n9062) );
  BUFx3_ASAP7_75t_R register___U13585 ( .A(register__n10219), .Y(register__n9063) );
  BUFx4f_ASAP7_75t_R register___U13586 ( .A(register__n6044), .Y(register__n9064) );
  BUFx12f_ASAP7_75t_R register___U13587 ( .A(register__n6045), .Y(register__n9810) );
  BUFx6f_ASAP7_75t_R register___U13588 ( .A(register__n9064), .Y(register__n9811) );
  BUFx4f_ASAP7_75t_R register___U13589 ( .A(register__n8024), .Y(register__n9066) );
  BUFx2_ASAP7_75t_R register___U13590 ( .A(Reg_data[124]), .Y(register__n9067) );
  BUFx12f_ASAP7_75t_R register___U13591 ( .A(register__n10224), .Y(register__n9068) );
  BUFx12f_ASAP7_75t_R register___U13592 ( .A(register__n9068), .Y(register__n10223) );
  BUFx6f_ASAP7_75t_R register___U13593 ( .A(register__n9066), .Y(register__n10224) );
  BUFx3_ASAP7_75t_R register___U13594 ( .A(register__n9070), .Y(register__n9069) );
  BUFx2_ASAP7_75t_R register___U13595 ( .A(Reg_data[444]), .Y(register__n9070) );
  BUFx4f_ASAP7_75t_R register___U13596 ( .A(register__n6812), .Y(register__n9071) );
  BUFx2_ASAP7_75t_R register___U13597 ( .A(Reg_data[883]), .Y(register__n9072) );
  BUFx12f_ASAP7_75t_R register___U13598 ( .A(register__n9825), .Y(register__n9073) );
  BUFx12f_ASAP7_75t_R register___U13599 ( .A(register__n9073), .Y(register__n9824) );
  BUFx6f_ASAP7_75t_R register___U13600 ( .A(register__n9071), .Y(register__n9825) );
  BUFx3_ASAP7_75t_R register___U13601 ( .A(register__n9075), .Y(register__n9074) );
  BUFx2_ASAP7_75t_R register___U13602 ( .A(Reg_data[115]), .Y(register__n9075) );
  BUFx12f_ASAP7_75t_R register___U13603 ( .A(register__n8025), .Y(register__n9076) );
  BUFx12f_ASAP7_75t_R register___U13604 ( .A(register__n9076), .Y(register__n10235) );
  BUFx3_ASAP7_75t_R register___U13605 ( .A(register__net94981), .Y(register__net94980) );
  BUFx2_ASAP7_75t_R register___U13606 ( .A(Reg_data[106]), .Y(register__net94981) );
  BUFx12f_ASAP7_75t_R register___U13607 ( .A(register__net89210), .Y(register__net89209) );
  BUFx3_ASAP7_75t_R register___U13608 ( .A(register__n9078), .Y(register__n9077) );
  BUFx2_ASAP7_75t_R register___U13609 ( .A(Reg_data[887]), .Y(register__n9078) );
  BUFx12f_ASAP7_75t_R register___U13610 ( .A(register__n9833), .Y(register__n9079) );
  BUFx12f_ASAP7_75t_R register___U13611 ( .A(register__n9079), .Y(register__n9832) );
  BUFx3_ASAP7_75t_R register___U13612 ( .A(register__n9081), .Y(register__n9080) );
  BUFx2_ASAP7_75t_R register___U13613 ( .A(Reg_data[695]), .Y(register__n9081) );
  BUFx12f_ASAP7_75t_R register___U13614 ( .A(register__n10262), .Y(register__n9082) );
  BUFx12f_ASAP7_75t_R register___U13615 ( .A(register__n9082), .Y(register__n10261) );
  BUFx3_ASAP7_75t_R register___U13616 ( .A(register__n9084), .Y(register__n9083) );
  BUFx2_ASAP7_75t_R register___U13617 ( .A(Reg_data[923]), .Y(register__n9084) );
  BUFx12f_ASAP7_75t_R register___U13618 ( .A(register__n9841), .Y(register__n9085) );
  BUFx12f_ASAP7_75t_R register___U13619 ( .A(register__n9085), .Y(register__n9840) );
  BUFx3_ASAP7_75t_R register___U13620 ( .A(register__n9087), .Y(register__n9086) );
  BUFx2_ASAP7_75t_R register___U13621 ( .A(Reg_data[247]), .Y(register__n9087) );
  BUFx12f_ASAP7_75t_R register___U13622 ( .A(register__n10272), .Y(register__n9088) );
  BUFx12f_ASAP7_75t_R register___U13623 ( .A(register__n9088), .Y(register__n10271) );
  BUFx3_ASAP7_75t_R register___U13624 ( .A(register__n9090), .Y(register__n9089) );
  BUFx2_ASAP7_75t_R register___U13625 ( .A(Reg_data[105]), .Y(register__n9090) );
  BUFx12f_ASAP7_75t_R register___U13626 ( .A(register__n10276), .Y(register__n9091) );
  BUFx12f_ASAP7_75t_R register___U13627 ( .A(register__n9091), .Y(register__n10275) );
  BUFx3_ASAP7_75t_R register___U13628 ( .A(register__n9093), .Y(register__n9092) );
  BUFx2_ASAP7_75t_R register___U13629 ( .A(Reg_data[762]), .Y(register__n9093) );
  BUFx2_ASAP7_75t_R register___U13630 ( .A(register__n9851), .Y(register__n9094) );
  BUFx2_ASAP7_75t_R register___U13631 ( .A(register__n9851), .Y(register__n9095) );
  BUFx4f_ASAP7_75t_R register___U13632 ( .A(register__n9851), .Y(register__n9096) );
  BUFx3_ASAP7_75t_R register___U13633 ( .A(register__n9098), .Y(register__n9097) );
  BUFx2_ASAP7_75t_R register___U13634 ( .A(Reg_data[698]), .Y(register__n9098) );
  BUFx12f_ASAP7_75t_R register___U13635 ( .A(register__n10290), .Y(register__n9099) );
  BUFx4f_ASAP7_75t_R register___U13636 ( .A(register__n6532), .Y(register__n9100) );
  BUFx2_ASAP7_75t_R register___U13637 ( .A(Reg_data[730]), .Y(register__n9101) );
  BUFx12f_ASAP7_75t_R register___U13638 ( .A(register__n10292), .Y(register__n9102) );
  BUFx12f_ASAP7_75t_R register___U13639 ( .A(register__n9102), .Y(register__n10291) );
  BUFx6f_ASAP7_75t_R register___U13640 ( .A(register__n9100), .Y(register__n10292) );
  BUFx4f_ASAP7_75t_R register___U13641 ( .A(register__n7709), .Y(register__n9103) );
  BUFx2_ASAP7_75t_R register___U13642 ( .A(Reg_data[895]), .Y(register__n9104) );
  BUFx12f_ASAP7_75t_R register___U13643 ( .A(register__n9858), .Y(register__n9857) );
  BUFx6f_ASAP7_75t_R register___U13644 ( .A(register__n9103), .Y(register__n9858) );
  BUFx3_ASAP7_75t_R register___U13645 ( .A(register__n9106), .Y(register__n9105) );
  BUFx2_ASAP7_75t_R register___U13646 ( .A(Reg_data[378]), .Y(register__n9106) );
  BUFx12f_ASAP7_75t_R register___U13647 ( .A(register__n9868), .Y(register__n9107) );
  BUFx12f_ASAP7_75t_R register___U13648 ( .A(register__n9107), .Y(register__n9867) );
  BUFx3_ASAP7_75t_R register___U13649 ( .A(register__n9109), .Y(register__n9108) );
  BUFx2_ASAP7_75t_R register___U13650 ( .A(Reg_data[410]), .Y(register__n9109) );
  BUFx2_ASAP7_75t_R register___U13651 ( .A(register__n9869), .Y(register__n9110) );
  BUFx2_ASAP7_75t_R register___U13652 ( .A(register__n9869), .Y(register__n9111) );
  BUFx4f_ASAP7_75t_R register___U13653 ( .A(register__n9869), .Y(register__n9112) );
  BUFx3_ASAP7_75t_R register___U13654 ( .A(register__n9114), .Y(register__n9113) );
  BUFx2_ASAP7_75t_R register___U13655 ( .A(Reg_data[58]), .Y(register__n9114) );
  BUFx12f_ASAP7_75t_R register___U13656 ( .A(register__n10302), .Y(register__n9115) );
  BUFx12f_ASAP7_75t_R register___U13657 ( .A(register__n9115), .Y(register__n10301) );
  BUFx3_ASAP7_75t_R register___U13658 ( .A(register__n9117), .Y(register__n9116) );
  BUFx2_ASAP7_75t_R register___U13659 ( .A(Reg_data[122]), .Y(register__n9117) );
  BUFx12f_ASAP7_75t_R register___U13660 ( .A(register__n8026), .Y(register__n9118) );
  BUFx12f_ASAP7_75t_R register___U13661 ( .A(register__n9118), .Y(register__n10303) );
  BUFx3_ASAP7_75t_R register___U13662 ( .A(register__n9120), .Y(register__n9119) );
  BUFx2_ASAP7_75t_R register___U13663 ( .A(Reg_data[108]), .Y(register__n9120) );
  BUFx12f_ASAP7_75t_R register___U13664 ( .A(register__n10306), .Y(register__n9121) );
  BUFx12f_ASAP7_75t_R register___U13665 ( .A(register__n9121), .Y(register__n10305) );
  BUFx3_ASAP7_75t_R register___U13666 ( .A(register__n9123), .Y(register__n9122) );
  BUFx2_ASAP7_75t_R register___U13667 ( .A(Reg_data[369]), .Y(register__n9123) );
  BUFx12f_ASAP7_75t_R register___U13668 ( .A(register__n9884), .Y(register__n9124) );
  BUFx12f_ASAP7_75t_R register___U13669 ( .A(register__n9124), .Y(register__n9883) );
  BUFx3_ASAP7_75t_R register___U13670 ( .A(register__net94863), .Y(register__net94862) );
  BUFx2_ASAP7_75t_R register___U13671 ( .A(Reg_data[888]), .Y(register__net94863) );
  BUFx12f_ASAP7_75t_R register___U13672 ( .A(register__net104001), .Y(register__net90257) );
  BUFx3_ASAP7_75t_R register___U13673 ( .A(register__n9126), .Y(register__n9125) );
  BUFx2_ASAP7_75t_R register___U13674 ( .A(Reg_data[127]), .Y(register__n9126) );
  BUFx12f_ASAP7_75t_R register___U13675 ( .A(register__n10328), .Y(register__n9127) );
  BUFx12f_ASAP7_75t_R register___U13676 ( .A(register__n9127), .Y(register__n10327) );
  BUFx3_ASAP7_75t_R register___U13677 ( .A(register__n9129), .Y(register__n9128) );
  BUFx2_ASAP7_75t_R register___U13678 ( .A(Reg_data[223]), .Y(register__n9129) );
  BUFx4f_ASAP7_75t_R register___U13679 ( .A(register__n10329), .Y(register__n9130) );
  BUFx2_ASAP7_75t_R register___U13680 ( .A(register__n10329), .Y(register__n9131) );
  BUFx3_ASAP7_75t_R register___U13681 ( .A(register__n10329), .Y(register__n9132) );
  BUFx4f_ASAP7_75t_R register___U13682 ( .A(register__n7710), .Y(register__n9133) );
  BUFx2_ASAP7_75t_R register___U13683 ( .A(Reg_data[31]), .Y(register__n9134) );
  BUFx12f_ASAP7_75t_R register___U13684 ( .A(register__n9136), .Y(register__n9135) );
  BUFx12f_ASAP7_75t_R register___U13685 ( .A(register__n10416), .Y(register__n9136) );
  BUFx12f_ASAP7_75t_R register___U13686 ( .A(register__n9135), .Y(register__n10415) );
  BUFx6f_ASAP7_75t_R register___U13687 ( .A(register__n9133), .Y(register__n10416) );
  BUFx4f_ASAP7_75t_R register___U13688 ( .A(register__n7711), .Y(register__n9137) );
  BUFx2_ASAP7_75t_R register___U13689 ( .A(Reg_data[95]), .Y(register__n9138) );
  BUFx12f_ASAP7_75t_R register___U13690 ( .A(register__n9140), .Y(register__n9139) );
  BUFx12f_ASAP7_75t_R register___U13691 ( .A(register__n10418), .Y(register__n9140) );
  BUFx12f_ASAP7_75t_R register___U13692 ( .A(register__n9139), .Y(register__n10417) );
  BUFx6f_ASAP7_75t_R register___U13693 ( .A(register__n9137), .Y(register__n10418) );
  BUFx4f_ASAP7_75t_R register___U13694 ( .A(register__net103992), .Y(register__net94817) );
  BUFx2_ASAP7_75t_R register___U13695 ( .A(Reg_data[29]), .Y(register__net94818) );
  BUFx12f_ASAP7_75t_R register___U13696 ( .A(register__net103991), .Y(register__net88764) );
  BUFx6f_ASAP7_75t_R register___U13697 ( .A(register__net94817), .Y(register__net88765) );
  BUFx4f_ASAP7_75t_R register___U13698 ( .A(register__net103988), .Y(register__net94809) );
  BUFx12f_ASAP7_75t_R register___U13699 ( .A(register__net103987), .Y(register__net88760) );
  BUFx6f_ASAP7_75t_R register___U13700 ( .A(register__net94809), .Y(register__net88761) );
  BUFx3_ASAP7_75t_R register___U13701 ( .A(register__net94800), .Y(register__net94799) );
  BUFx2_ASAP7_75t_R register___U13702 ( .A(Reg_data[893]), .Y(register__net94800) );
  BUFx2_ASAP7_75t_R register___U13703 ( .A(register__net90221), .Y(register__net94801) );
  BUFx4f_ASAP7_75t_R register___U13704 ( .A(register__net90221), .Y(register__net94803) );
  BUFx3_ASAP7_75t_R register___U13705 ( .A(register__net94796), .Y(register__net94795) );
  BUFx2_ASAP7_75t_R register___U13706 ( .A(Reg_data[669]), .Y(register__net94796) );
  BUFx3_ASAP7_75t_R register___U13707 ( .A(register__net94786), .Y(register__net94785) );
  BUFx2_ASAP7_75t_R register___U13708 ( .A(Reg_data[733]), .Y(register__net94786) );
  BUFx4f_ASAP7_75t_R register___U13709 ( .A(register__net88997), .Y(register__net94787) );
  BUFx3_ASAP7_75t_R register___U13710 ( .A(register__net88997), .Y(register__net94789) );
  BUFx4f_ASAP7_75t_R register___U13711 ( .A(register__net103985), .Y(register__net94775) );
  BUFx2_ASAP7_75t_R register___U13712 ( .A(Reg_data[797]), .Y(register__net94776) );
  BUFx12f_ASAP7_75t_R register___U13713 ( .A(register__net94778), .Y(register__net88756) );
  BUFx12f_ASAP7_75t_R register___U13714 ( .A(register__net88757), .Y(register__net94778) );
  BUFx6f_ASAP7_75t_R register___U13715 ( .A(register__net94775), .Y(register__net88757) );
  BUFx4f_ASAP7_75t_R register___U13716 ( .A(register__net103982), .Y(register__net94767) );
  BUFx2_ASAP7_75t_R register___U13717 ( .A(Reg_data[861]), .Y(register__net94768) );
  BUFx12f_ASAP7_75t_R register___U13718 ( .A(register__net103981), .Y(register__net88752) );
  BUFx6f_ASAP7_75t_R register___U13719 ( .A(register__net94767), .Y(register__net88753) );
  BUFx3_ASAP7_75t_R register___U13720 ( .A(register__n9142), .Y(register__n9141) );
  BUFx2_ASAP7_75t_R register___U13721 ( .A(Reg_data[892]), .Y(register__n9142) );
  BUFx12f_ASAP7_75t_R register___U13722 ( .A(register__n9898), .Y(register__n9897) );
  BUFx3_ASAP7_75t_R register___U13723 ( .A(register__n9144), .Y(register__n9143) );
  BUFx2_ASAP7_75t_R register___U13724 ( .A(Reg_data[668]), .Y(register__n9144) );
  BUFx12f_ASAP7_75t_R register___U13725 ( .A(register__n6282), .Y(register__n10335) );
  BUFx3_ASAP7_75t_R register___U13726 ( .A(register__n9146), .Y(register__n9145) );
  BUFx2_ASAP7_75t_R register___U13727 ( .A(Reg_data[478]), .Y(register__n9146) );
  BUFx12f_ASAP7_75t_R register___U13728 ( .A(register__n9910), .Y(register__n9147) );
  BUFx12f_ASAP7_75t_R register___U13729 ( .A(register__n9147), .Y(register__n9909) );
  BUFx6f_ASAP7_75t_R register___U13730 ( .A(register__n4866), .Y(register__n12036) );
  BUFx6f_ASAP7_75t_R register___U13731 ( .A(register__n3837), .Y(register__n12038) );
  BUFx4f_ASAP7_75t_R register___U13732 ( .A(register__n4866), .Y(register__n12039) );
  BUFx12f_ASAP7_75t_R register___U13733 ( .A(register__n4865), .Y(register__n12049) );
  INVx1_ASAP7_75t_R register___U13734 ( .A(register__n5416), .Y(register__n9149) );
  INVx1_ASAP7_75t_R register___U13735 ( .A(register__n5418), .Y(register__n9150) );
  INVx1_ASAP7_75t_R register___U13736 ( .A(register__n5420), .Y(register__n9151) );
  INVx1_ASAP7_75t_R register___U13737 ( .A(register__n4991), .Y(register__n9152) );
  INVx1_ASAP7_75t_R register___U13738 ( .A(register__n5066), .Y(register__n9153) );
  BUFx6f_ASAP7_75t_R register___U13739 ( .A(register__n4748), .Y(register__n12178) );
  INVx3_ASAP7_75t_R register___U13740 ( .A(register__net99033), .Y(register__net94613) );
  INVx3_ASAP7_75t_R register___U13741 ( .A(register__n11623), .Y(register__n9159) );
  INVx2_ASAP7_75t_R register___U13742 ( .A(register__n11181), .Y(register__n9160) );
  BUFx2_ASAP7_75t_R register___U13743 ( .A(Reg_data[593]), .Y(register__n10845) );
  INVx2_ASAP7_75t_R register___U13744 ( .A(register__n6778), .Y(register__n9161) );
  OA22x2_ASAP7_75t_R register___U13745 ( .A1(register__n12323), .A2(register__n7327), .B1(register__n5190), .B2(register__n3505), 
        .Y(register__n12561) );
  INVx1_ASAP7_75t_R register___U13746 ( .A(register__n12561), .Y(register__n9162) );
  OA22x2_ASAP7_75t_R register___U13747 ( .A1(register__net64944), .A2(register__n7327), .B1(register__n9589), .B2(register__n4818), .Y(register__n12574) );
  INVx1_ASAP7_75t_R register___U13748 ( .A(register__n12574), .Y(register__n9163) );
  OA22x2_ASAP7_75t_R register___U13749 ( .A1(register__net64664), .A2(register__n7327), .B1(register__n7801), .B2(register__n3947), .Y(register__n12571) );
  OA22x2_ASAP7_75t_R register___U13750 ( .A1(register__n12124), .A2(register__n7327), .B1(register__n9816), .B2(register__n11912), 
        .Y(register__n12567) );
  INVx4_ASAP7_75t_R register___U13751 ( .A(register__n12138), .Y(register__n12124) );
  OA22x2_ASAP7_75t_R register___U13752 ( .A1(register__n12407), .A2(register__n7327), .B1(register__n9855), .B2(register__n89), 
        .Y(register__n12557) );
  INVx1_ASAP7_75t_R register___U13753 ( .A(register__n12557), .Y(register__n9166) );
  OA22x2_ASAP7_75t_R register___U13754 ( .A1(register__n12093), .A2(register__n7327), .B1(register__n7554), .B2(register__n11835), 
        .Y(register__n12569) );
  OA22x2_ASAP7_75t_R register___U13755 ( .A1(register__net63264), .A2(register__n7327), .B1(register__net90249), .B2(
        n3472), .Y(register__n12559) );
  INVx1_ASAP7_75t_R register___U13756 ( .A(register__n12559), .Y(register__n9167) );
  AO22x1_ASAP7_75t_R register___U13757 ( .A1(register__n8795), .A2(register__C6423_net61318), .B1(register__n8349), 
        .B2(register__n1449), .Y(register__n11186) );
  INVx1_ASAP7_75t_R register___U13758 ( .A(register__n4734), .Y(register__n9168) );
  BUFx6f_ASAP7_75t_R register___U13759 ( .A(register__n12012), .Y(register__n12000) );
  BUFx12f_ASAP7_75t_R register___U13760 ( .A(register__n12017), .Y(register__n12016) );
  BUFx6f_ASAP7_75t_R register___U13761 ( .A(register__n4746), .Y(register__n12307) );
  BUFx6f_ASAP7_75t_R register___U13762 ( .A(register__net121483), .Y(register__net62866) );
  BUFx6f_ASAP7_75t_R register___U13763 ( .A(register__net62848), .Y(register__net62876) );
  BUFx6f_ASAP7_75t_R register___U13764 ( .A(register__net121484), .Y(register__net62870) );
  BUFx6f_ASAP7_75t_R register___U13765 ( .A(register__net140665), .Y(register__net62878) );
  OA22x2_ASAP7_75t_R register___U13766 ( .A1(register__n11963), .A2(register__n11915), .B1(register__n5199), .B2(register__n3506), 
        .Y(register__n12577) );
  INVx1_ASAP7_75t_R register___U13767 ( .A(register__n5392), .Y(register__n9171) );
  INVx1_ASAP7_75t_R register___U13768 ( .A(register__n2991), .Y(register__n9172) );
  INVx1_ASAP7_75t_R register___U13769 ( .A(register__n2993), .Y(register__n9173) );
  INVx1_ASAP7_75t_R register___U13770 ( .A(register__n2995), .Y(register__n9174) );
  AO22x1_ASAP7_75t_R register___U13771 ( .A1(register__net104596), .A2(register__C6423_net61318), .B1(
        net89861), .B2(register__n1446), .Y(register__n11268) );
  AO22x1_ASAP7_75t_R register___U13772 ( .A1(register__net96915), .A2(register__n156), .B1(register__net89013), .B2(
        n281), .Y(register__n11096) );
  INVx1_ASAP7_75t_R register___U13773 ( .A(register__n11096), .Y(register__n9181) );
  OA22x2_ASAP7_75t_R register___U13774 ( .A1(register__n3253), .A2(register__n111), .B1(register__n9549), .B2(register__n1662), 
        .Y(register__n12651) );
  OA22x2_ASAP7_75t_R register___U13775 ( .A1(register__n11816), .A2(register__n12235), .B1(register__n9571), .B2(register__n1598), 
        .Y(register__n12702) );
  OA22x2_ASAP7_75t_R register___U13776 ( .A1(register__n12434), .A2(register__n7327), .B1(register__n9901), .B2(register__n5171), 
        .Y(register__n12556) );
  INVx1_ASAP7_75t_R register___U13777 ( .A(register__n4601), .Y(register__n9185) );
  OR3x1_ASAP7_75t_R register___U13778 ( .A(register__n7362), .B(register__n9188), .C(register__n9187), .Y(register__n10570) );
  OA22x2_ASAP7_75t_R register___U13779 ( .A1(register__n420), .A2(register__n6486), .B1(register__n801), .B2(register__n11202), 
        .Y(register__n10573) );
  INVx1_ASAP7_75t_R register___U13780 ( .A(register__n7358), .Y(register__n9187) );
  OA22x2_ASAP7_75t_R register___U13781 ( .A1(register__n66), .A2(register__n11203), .B1(register__n1691), .B2(register__n7692), 
        .Y(register__n10572) );
  OA222x2_ASAP7_75t_R register___U13782 ( .A1(register__n2002), .A2(register__n11204), .B1(register__n1997), .B2(register__n11205), .C1(register__net112580), .C2(register__n11206), .Y(register__n10571) );
  OR3x1_ASAP7_75t_R register___U13783 ( .A(register__n533), .B(register__n9191), .C(register__n9190), .Y(register__n11099) );
  OA22x2_ASAP7_75t_R register___U13784 ( .A1(register__n420), .A2(register__register__n8005), .B1(register__n800), .B2(register__n11686), 
        .Y(register__n11102) );
  INVx1_ASAP7_75t_R register___U13785 ( .A(register__n7698), .Y(register__n9190) );
  OA22x2_ASAP7_75t_R register___U13786 ( .A1(register__net107674), .A2(register__n7099), .B1(register__n1691), .B2(
        n7345), .Y(register__n11101) );
  OA222x2_ASAP7_75t_R register___U13787 ( .A1(register__n2002), .A2(register__n6475), .B1(register__net130666), .B2(
        n11107), .C1(register__net112580), .C2(register__n6211), .Y(register__n11100) );
  OR3x1_ASAP7_75t_R register___U13788 ( .A(register__n9194), .B(register__n9193), .C(register__n9192), .Y(register__n11681) );
  OA22x2_ASAP7_75t_R register___U13789 ( .A1(register__net131654), .A2(register__n6491), .B1(register__net130175), .B2(
        n8008), .Y(register__n11684) );
  INVx1_ASAP7_75t_R register___U13790 ( .A(register__n5476), .Y(register__n9192) );
  OA22x2_ASAP7_75t_R register___U13791 ( .A1(register__n713), .A2(register__n11104), .B1(register__net149934), .B2(
        n11105), .Y(register__n11683) );
  INVx1_ASAP7_75t_R register___U13792 ( .A(register__n5478), .Y(register__n9193) );
  OA222x2_ASAP7_75t_R register___U13793 ( .A1(register__n1987), .A2(register__n11106), .B1(register__n1995), .B2(register__n11687), .C1(register__n1800), .C2(register__n11108), .Y(register__n11682) );
  OR3x1_ASAP7_75t_R register___U13794 ( .A(register__n9196), .B(register__n258), .C(register__n9195), .Y(register__n10951) );
  OA22x2_ASAP7_75t_R register___U13795 ( .A1(register__n420), .A2(register__n6487), .B1(register__n800), .B2(register__n6777), 
        .Y(register__n10954) );
  INVx1_ASAP7_75t_R register___U13796 ( .A(register__n5455), .Y(register__n9195) );
  OA22x2_ASAP7_75t_R register___U13797 ( .A1(register__net107674), .A2(register__n11567), .B1(register__n1691), .B2(
        n7342), .Y(register__n10953) );
  OA222x2_ASAP7_75t_R register___U13798 ( .A1(register__n2002), .A2(register__n6218), .B1(register__n817), .B2(register__n5953), 
        .C1(register__net112580), .C2(register__n5725), .Y(register__n10952) );
  INVx1_ASAP7_75t_R register___U13799 ( .A(register__n10952), .Y(register__n9196) );
  OA22x2_ASAP7_75t_R register___U13800 ( .A1(register__n420), .A2(register__net111143), .B1(register__n800), .B2(
        net104283), .Y(register__n10720) );
  INVx1_ASAP7_75t_R register___U13801 ( .A(register__n4829), .Y(register__n9197) );
  OA22x2_ASAP7_75t_R register___U13802 ( .A1(register__net107674), .A2(register__C6423_net60775), .B1(register__n1691), 
        .B2(register__net105518), .Y(register__n10719) );
  INVx1_ASAP7_75t_R register___U13803 ( .A(register__n4831), .Y(register__n9198) );
  OA222x2_ASAP7_75t_R register___U13804 ( .A1(register__n2080), .A2(register__C6423_net60777), .B1(register__n1997), 
        .B2(register__C6422_net59860), .C1(register__C6422_net69812), .C2(register__net107836), .Y(register__n10718)
         );
  INVx1_ASAP7_75t_R register___U13805 ( .A(register__n4833), .Y(register__n9199) );
  OR3x1_ASAP7_75t_R register___U13806 ( .A(register__n5636), .B(register__n9201), .C(register__n9200), .Y(register__n11602) );
  OA22x2_ASAP7_75t_R register___U13807 ( .A1(register__net131654), .A2(register__net99209), .B1(register__net130175), 
        .B2(register__net105510), .Y(register__n11605) );
  INVx1_ASAP7_75t_R register___U13808 ( .A(register__n5632), .Y(register__n9200) );
  OA22x2_ASAP7_75t_R register___U13809 ( .A1(register__n712), .A2(register__net111131), .B1(register__n353), .B2(
        net108759), .Y(register__n11604) );
  INVx1_ASAP7_75t_R register___U13810 ( .A(register__n5634), .Y(register__n9201) );
  OA222x2_ASAP7_75t_R register___U13811 ( .A1(register__n1987), .A2(register__C6423_net61115), .B1(register__n1995), 
        .B2(register__C6423_net61116), .C1(register__n1800), .C2(register__net103314), .Y(register__n11603) );
  OR3x1_ASAP7_75t_R register___U13812 ( .A(register__n5488), .B(register__n9204), .C(register__n9203), .Y(register__n11037) );
  OA22x2_ASAP7_75t_R register___U13813 ( .A1(register__n419), .A2(register__n7347), .B1(register__n802), .B2(register__n11644), 
        .Y(register__n11040) );
  INVx1_ASAP7_75t_R register___U13814 ( .A(register__n5482), .Y(register__n9203) );
  OA22x2_ASAP7_75t_R register___U13815 ( .A1(register__n66), .A2(register__n11645), .B1(register__n1691), .B2(register__n11042), 
        .Y(register__n11039) );
  INVx1_ASAP7_75t_R register___U13816 ( .A(register__n5484), .Y(register__n9204) );
  OA222x2_ASAP7_75t_R register___U13817 ( .A1(register__n2002), .A2(register__n7090), .B1(register__n817), .B2(
        C6423_net61194), .C1(register__net112580), .C2(register__net103310), .Y(register__n11038) );
  INVx1_ASAP7_75t_R register___U13818 ( .A(register__n5486), .Y(register__n9205) );
  OA22x2_ASAP7_75t_R register___U13819 ( .A1(register__n1965), .A2(register__n6492), .B1(register__net130175), .B2(
        n8590), .Y(register__n11370) );
  OA22x2_ASAP7_75t_R register___U13820 ( .A1(register__n713), .A2(register__n10741), .B1(register__n353), .B2(register__n7109), 
        .Y(register__n11369) );
  INVx1_ASAP7_75t_R register___U13821 ( .A(register__n6023), .Y(register__n9207) );
  OA222x2_ASAP7_75t_R register___U13822 ( .A1(register__n1987), .A2(register__n5731), .B1(register__n1995), .B2(register__n10743), 
        .C1(register__n1800), .C2(register__n7578), .Y(register__n11368) );
  BUFx3_ASAP7_75t_R register___U13823 ( .A(register__n8373), .Y(register__n9210) );
  BUFx3_ASAP7_75t_R register___U13824 ( .A(register__net98827), .Y(register__net94161) );
  OA22x2_ASAP7_75t_R register___U13825 ( .A1(register__n2013), .A2(register__n8002), .B1(register__net130175), .B2(
        n6769), .Y(register__n11200) );
  INVx1_ASAP7_75t_R register___U13826 ( .A(register__n11200), .Y(register__n9219) );
  OA22x2_ASAP7_75t_R register___U13827 ( .A1(register__n711), .A2(register__n7690), .B1(register__n1113), .B2(register__n10575), 
        .Y(register__n11199) );
  INVx1_ASAP7_75t_R register___U13828 ( .A(register__n5334), .Y(register__n9221) );
  OA22x2_ASAP7_75t_R register___U13829 ( .A1(register__n1965), .A2(register__n6770), .B1(register__net130175), .B2(
        n10530), .Y(register__n11159) );
  INVx1_ASAP7_75t_R register___U13830 ( .A(register__n6001), .Y(register__n9222) );
  OA22x2_ASAP7_75t_R register___U13831 ( .A1(register__n713), .A2(register__n7869), .B1(register__n10531), .B2(register__n353), 
        .Y(register__n11158) );
  INVx1_ASAP7_75t_R register___U13832 ( .A(register__n6006), .Y(register__n9224) );
  OR3x1_ASAP7_75t_R register___U13833 ( .A(register__n9227), .B(register__n9226), .C(register__n9225), .Y(register__n10782) );
  OA22x2_ASAP7_75t_R register___U13834 ( .A1(register__n66), .A2(register__n10787), .B1(register__n1691), .B2(register__n7585), 
        .Y(register__n10784) );
  OA222x2_ASAP7_75t_R register___U13835 ( .A1(register__n2080), .A2(register__n6478), .B1(register__n1117), .B2(register__n11415), 
        .C1(register__net112580), .C2(register__n5954), .Y(register__n10783) );
  INVx1_ASAP7_75t_R register___U13836 ( .A(register__n5474), .Y(register__n9227) );
  OR3x1_ASAP7_75t_R register___U13837 ( .A(register__n9230), .B(register__n9229), .C(register__n9228), .Y(register__n10862) );
  OA22x2_ASAP7_75t_R register___U13838 ( .A1(register__n420), .A2(register__n7096), .B1(register__n800), .B2(register__n6772), 
        .Y(register__n10865) );
  INVx1_ASAP7_75t_R register___U13839 ( .A(register__n4938), .Y(register__n9228) );
  OA22x2_ASAP7_75t_R register___U13840 ( .A1(register__net107674), .A2(register__n7870), .B1(register__n1691), .B2(
        n6481), .Y(register__n10864) );
  INVx1_ASAP7_75t_R register___U13841 ( .A(register__n4940), .Y(register__n9229) );
  OA222x2_ASAP7_75t_R register___U13842 ( .A1(register__n2002), .A2(register__n6216), .B1(register__n817), .B2(register__n7579), 
        .C1(register__net112580), .C2(register__n11482), .Y(register__n10863) );
  INVx1_ASAP7_75t_R register___U13843 ( .A(register__n4942), .Y(register__n9230) );
  OA22x2_ASAP7_75t_R register___U13844 ( .A1(register__n66), .A2(register__n11350), .B1(register__n1691), .B2(register__n7582), 
        .Y(register__n10681) );
  OA222x2_ASAP7_75t_R register___U13845 ( .A1(register__n2080), .A2(register__n6222), .B1(register__n817), .B2(register__n11352), 
        .C1(register__net112580), .C2(register__n11353), .Y(register__n10680) );
  OR3x1_ASAP7_75t_R register___U13846 ( .A(register__n5446), .B(register__n9235), .C(register__n9233), .Y(register__n11281) );
  OA22x2_ASAP7_75t_R register___U13847 ( .A1(register__net131654), .A2(register__net106698), .B1(register__net130175), 
        .B2(register__C6422_net59726), .Y(register__n11284) );
  INVx1_ASAP7_75t_R register___U13848 ( .A(register__n5444), .Y(register__n9233) );
  OA222x2_ASAP7_75t_R register___U13849 ( .A1(register__n1987), .A2(register__C6422_net59729), .B1(register__n1995), 
        .B2(register__C6422_net59730), .C1(register__n1800), .C2(register__C6422_net59731), .Y(register__n11282) );
  INVx1_ASAP7_75t_R register___U13850 ( .A(register__n11282), .Y(register__n9234) );
  OA22x2_ASAP7_75t_R register___U13851 ( .A1(register__n712), .A2(register__net108801), .B1(register__n407), .B2(
        net100833), .Y(register__n11283) );
  INVx1_ASAP7_75t_R register___U13852 ( .A(register__n5447), .Y(register__n9235) );
  OR3x1_ASAP7_75t_R register___U13853 ( .A(register__n7369), .B(register__n9237), .C(register__n9236), .Y(register__n11659) );
  OA22x2_ASAP7_75t_R register___U13854 ( .A1(register__n711), .A2(register__n11061), .B1(register__n353), .B2(register__n11062), 
        .Y(register__n11661) );
  INVx1_ASAP7_75t_R register___U13855 ( .A(register__n7365), .Y(register__n9237) );
  OA222x2_ASAP7_75t_R register___U13856 ( .A1(register__net127626), .A2(register__n11063), .B1(register__n1995), .B2(
        n11665), .C1(register__n1800), .C2(register__n11065), .Y(register__n11660) );
  OR3x1_ASAP7_75t_R register___U13857 ( .A(register__n6013), .B(register__n9240), .C(register__n9239), .Y(register__n11496) );
  OA22x2_ASAP7_75t_R register___U13858 ( .A1(register__C6423_net68482), .A2(register__n10890), .B1(register__net130175), 
        .B2(register__n8591), .Y(register__n11499) );
  OA22x2_ASAP7_75t_R register___U13859 ( .A1(register__n711), .A2(register__n7105), .B1(register__net149933), .B2(register__n7583), .Y(register__n11498) );
  INVx1_ASAP7_75t_R register___U13860 ( .A(register__n6011), .Y(register__n9240) );
  OR3x1_ASAP7_75t_R register___U13861 ( .A(register__n5994), .B(register__n9243), .C(register__n9242), .Y(register__n11543) );
  INVx1_ASAP7_75t_R register___U13862 ( .A(register__n5992), .Y(register__n9242) );
  OA22x2_ASAP7_75t_R register___U13863 ( .A1(register__n713), .A2(register__n10935), .B1(register__n353), .B2(register__n10936), 
        .Y(register__n11545) );
  INVx1_ASAP7_75t_R register___U13864 ( .A(register__n11545), .Y(register__n9243) );
  OA222x2_ASAP7_75t_R register___U13865 ( .A1(register__n1987), .A2(register__n6474), .B1(register__n1995), .B2(register__n7581), 
        .C1(register__n1800), .C2(register__n7866), .Y(register__n11544) );
  BUFx6f_ASAP7_75t_R register___U13866 ( .A(register__n9245), .Y(register__n9244) );
  BUFx4f_ASAP7_75t_R register___U13867 ( .A(register__n8471), .Y(register__n9245) );
  BUFx6f_ASAP7_75t_R register___U13868 ( .A(register__n9247), .Y(register__n9246) );
  BUFx4f_ASAP7_75t_R register___U13869 ( .A(register__n6107), .Y(register__n9247) );
  BUFx4f_ASAP7_75t_R register___U13870 ( .A(register__net116146), .Y(register__net93853) );
  BUFx6f_ASAP7_75t_R register___U13871 ( .A(register__n9249), .Y(register__n9248) );
  BUFx4f_ASAP7_75t_R register___U13872 ( .A(register__n5845), .Y(register__n9249) );
  BUFx6f_ASAP7_75t_R register___U13873 ( .A(register__n9251), .Y(register__n9250) );
  BUFx4f_ASAP7_75t_R register___U13874 ( .A(register__n6831), .Y(register__n9251) );
  BUFx6f_ASAP7_75t_R register___U13875 ( .A(register__n9253), .Y(register__n9252) );
  BUFx4f_ASAP7_75t_R register___U13876 ( .A(register__n6303), .Y(register__n9253) );
  BUFx4f_ASAP7_75t_R register___U13877 ( .A(register__net116142), .Y(register__net93837) );
  BUFx6f_ASAP7_75t_R register___U13878 ( .A(register__n9255), .Y(register__n9254) );
  BUFx4f_ASAP7_75t_R register___U13879 ( .A(register__n5357), .Y(register__n9255) );
  BUFx6f_ASAP7_75t_R register___U13880 ( .A(register__n9257), .Y(register__n9256) );
  BUFx4f_ASAP7_75t_R register___U13881 ( .A(register__n7734), .Y(register__n9257) );
  BUFx6f_ASAP7_75t_R register___U13882 ( .A(register__n9259), .Y(register__n9258) );
  BUFx4f_ASAP7_75t_R register___U13883 ( .A(register__n6340), .Y(register__n9259) );
  BUFx6f_ASAP7_75t_R register___U13884 ( .A(register__n9261), .Y(register__n9260) );
  BUFx4f_ASAP7_75t_R register___U13885 ( .A(register__n7177), .Y(register__n9261) );
  BUFx4f_ASAP7_75t_R register___U13886 ( .A(register__net114208), .Y(register__net93817) );
  BUFx6f_ASAP7_75t_R register___U13887 ( .A(register__n9263), .Y(register__n9262) );
  BUFx4f_ASAP7_75t_R register___U13888 ( .A(register__n6344), .Y(register__n9263) );
  BUFx6f_ASAP7_75t_R register___U13889 ( .A(register__n9265), .Y(register__n9264) );
  BUFx4f_ASAP7_75t_R register___U13890 ( .A(register__n6094), .Y(register__n9265) );
  BUFx4f_ASAP7_75t_R register___U13891 ( .A(register__net114200), .Y(register__net93805) );
  BUFx6f_ASAP7_75t_R register___U13892 ( .A(register__n9267), .Y(register__n9266) );
  BUFx4f_ASAP7_75t_R register___U13893 ( .A(register__n6597), .Y(register__n9267) );
  BUFx4f_ASAP7_75t_R register___U13894 ( .A(register__net112419), .Y(register__net93797) );
  BUFx4f_ASAP7_75t_R register___U13895 ( .A(register__net116044), .Y(register__net93793) );
  BUFx6f_ASAP7_75t_R register___U13896 ( .A(register__n9269), .Y(register__n9268) );
  BUFx4f_ASAP7_75t_R register___U13897 ( .A(register__n5528), .Y(register__n9269) );
  BUFx6f_ASAP7_75t_R register___U13898 ( .A(register__n9271), .Y(register__n9270) );
  BUFx4f_ASAP7_75t_R register___U13899 ( .A(register__n6105), .Y(register__n9271) );
  BUFx6f_ASAP7_75t_R register___U13900 ( .A(register__n9273), .Y(register__n9272) );
  BUFx4f_ASAP7_75t_R register___U13901 ( .A(register__n6358), .Y(register__n9273) );
  BUFx6f_ASAP7_75t_R register___U13902 ( .A(register__n9275), .Y(register__n9274) );
  BUFx4f_ASAP7_75t_R register___U13903 ( .A(register__n8098), .Y(register__n9275) );
  BUFx6f_ASAP7_75t_R register___U13904 ( .A(register__n9277), .Y(register__n9276) );
  BUFx4f_ASAP7_75t_R register___U13905 ( .A(register__n6894), .Y(register__n9277) );
  BUFx6f_ASAP7_75t_R register___U13906 ( .A(register__n9279), .Y(register__n9278) );
  BUFx4f_ASAP7_75t_R register___U13907 ( .A(register__n6899), .Y(register__n9279) );
  BUFx6f_ASAP7_75t_R register___U13908 ( .A(register__n9281), .Y(register__n9280) );
  BUFx4f_ASAP7_75t_R register___U13909 ( .A(register__n6901), .Y(register__n9281) );
  BUFx6f_ASAP7_75t_R register___U13910 ( .A(register__n9283), .Y(register__n9282) );
  BUFx4f_ASAP7_75t_R register___U13911 ( .A(register__n6613), .Y(register__n9283) );
  BUFx6f_ASAP7_75t_R register___U13912 ( .A(register__n9285), .Y(register__n9284) );
  BUFx4f_ASAP7_75t_R register___U13913 ( .A(register__n6615), .Y(register__n9285) );
  BUFx4f_ASAP7_75t_R register___U13914 ( .A(register__net110086), .Y(register__net93753) );
  BUFx6f_ASAP7_75t_R register___U13915 ( .A(register__n9287), .Y(register__n9286) );
  BUFx4f_ASAP7_75t_R register___U13916 ( .A(register__n6371), .Y(register__n9287) );
  BUFx6f_ASAP7_75t_R register___U13917 ( .A(register__n9289), .Y(register__n9288) );
  BUFx4f_ASAP7_75t_R register___U13918 ( .A(register__n6617), .Y(register__n9289) );
  BUFx4f_ASAP7_75t_R register___U13919 ( .A(register__net110082), .Y(register__net93741) );
  BUFx4f_ASAP7_75t_R register___U13920 ( .A(register__net110078), .Y(register__net93737) );
  BUFx6f_ASAP7_75t_R register___U13921 ( .A(register__n9291), .Y(register__n9290) );
  BUFx4f_ASAP7_75t_R register___U13922 ( .A(register__n6903), .Y(register__n9291) );
  BUFx6f_ASAP7_75t_R register___U13923 ( .A(register__n9293), .Y(register__n9292) );
  BUFx4f_ASAP7_75t_R register___U13924 ( .A(register__n6905), .Y(register__n9293) );
  BUFx6f_ASAP7_75t_R register___U13925 ( .A(register__n9295), .Y(register__n9294) );
  BUFx4f_ASAP7_75t_R register___U13926 ( .A(register__n6907), .Y(register__n9295) );
  BUFx4f_ASAP7_75t_R register___U13927 ( .A(register__net114119), .Y(register__net93717) );
  BUFx4f_ASAP7_75t_R register___U13928 ( .A(register__net112335), .Y(register__net93713) );
  BUFx4f_ASAP7_75t_R register___U13929 ( .A(register__n8481), .Y(register__n9298) );
  BUFx6f_ASAP7_75t_R register___U13930 ( .A(register__n9300), .Y(register__n9299) );
  BUFx4f_ASAP7_75t_R register___U13931 ( .A(register__n8145), .Y(register__n9300) );
  BUFx6f_ASAP7_75t_R register___U13932 ( .A(register__n9302), .Y(register__n9301) );
  BUFx4f_ASAP7_75t_R register___U13933 ( .A(register__n7523), .Y(register__n9302) );
  BUFx6f_ASAP7_75t_R register___U13934 ( .A(register__n9304), .Y(register__n9303) );
  BUFx4f_ASAP7_75t_R register___U13935 ( .A(register__n6640), .Y(register__n9304) );
  BUFx6f_ASAP7_75t_R register___U13936 ( .A(register__n9306), .Y(register__n9305) );
  BUFx4f_ASAP7_75t_R register___U13937 ( .A(register__n6953), .Y(register__n9306) );
  BUFx6f_ASAP7_75t_R register___U13938 ( .A(register__n9308), .Y(register__n9307) );
  BUFx4f_ASAP7_75t_R register___U13939 ( .A(register__n6652), .Y(register__n9308) );
  BUFx6f_ASAP7_75t_R register___U13940 ( .A(register__n9310), .Y(register__n9309) );
  BUFx4f_ASAP7_75t_R register___U13941 ( .A(register__n8512), .Y(register__n9310) );
  BUFx6f_ASAP7_75t_R register___U13942 ( .A(register__n9312), .Y(register__n9311) );
  BUFx4f_ASAP7_75t_R register___U13943 ( .A(register__n6962), .Y(register__n9312) );
  BUFx6f_ASAP7_75t_R register___U13944 ( .A(register__n9314), .Y(register__n9313) );
  BUFx4f_ASAP7_75t_R register___U13945 ( .A(register__n6666), .Y(register__n9314) );
  BUFx4f_ASAP7_75t_R register___U13946 ( .A(register__net107856), .Y(register__net93673) );
  BUFx6f_ASAP7_75t_R register___U13947 ( .A(register__n9316), .Y(register__n9315) );
  BUFx4f_ASAP7_75t_R register___U13948 ( .A(register__n6976), .Y(register__n9316) );
  BUFx6f_ASAP7_75t_R register___U13949 ( .A(register__n9318), .Y(register__n9317) );
  BUFx4f_ASAP7_75t_R register___U13950 ( .A(register__n6978), .Y(register__n9318) );
  BUFx6f_ASAP7_75t_R register___U13951 ( .A(register__n9320), .Y(register__n9319) );
  BUFx4f_ASAP7_75t_R register___U13952 ( .A(register__n8461), .Y(register__n9320) );
  BUFx6f_ASAP7_75t_R register___U13953 ( .A(register__n9322), .Y(register__n9321) );
  BUFx4f_ASAP7_75t_R register___U13954 ( .A(register__n5675), .Y(register__n9322) );
  BUFx4f_ASAP7_75t_R register___U13955 ( .A(register__net116040), .Y(register__net93639) );
  BUFx6f_ASAP7_75t_R register___U13956 ( .A(register__n9324), .Y(register__n9323) );
  BUFx4f_ASAP7_75t_R register___U13957 ( .A(register__n7157), .Y(register__n9324) );
  BUFx6f_ASAP7_75t_R register___U13958 ( .A(register__n9326), .Y(register__n9325) );
  BUFx4f_ASAP7_75t_R register___U13959 ( .A(register__n6315), .Y(register__n9326) );
  BUFx6f_ASAP7_75t_R register___U13960 ( .A(register__n9328), .Y(register__n9327) );
  BUFx4f_ASAP7_75t_R register___U13961 ( .A(register__n7509), .Y(register__n9328) );
  BUFx6f_ASAP7_75t_R register___U13962 ( .A(register__net93577), .Y(register__net93576) );
  BUFx4f_ASAP7_75t_R register___U13963 ( .A(register__net98494), .Y(register__net93577) );
  BUFx6f_ASAP7_75t_R register___U13964 ( .A(register__n9330), .Y(register__n9329) );
  BUFx4f_ASAP7_75t_R register___U13965 ( .A(register__n5851), .Y(register__n9330) );
  BUFx4f_ASAP7_75t_R register___U13966 ( .A(register__net114310), .Y(register__net93508) );
  BUFx6f_ASAP7_75t_R register___U13967 ( .A(register__n9332), .Y(register__n9331) );
  BUFx4f_ASAP7_75t_R register___U13968 ( .A(register__n6858), .Y(register__n9332) );
  BUFx6f_ASAP7_75t_R register___U13969 ( .A(register__n9336), .Y(register__n9335) );
  BUFx4f_ASAP7_75t_R register___U13970 ( .A(register__n8052), .Y(register__n9336) );
  BUFx6f_ASAP7_75t_R register___U13971 ( .A(register__n9338), .Y(register__n9337) );
  BUFx4f_ASAP7_75t_R register___U13972 ( .A(register__n6342), .Y(register__n9338) );
  BUFx6f_ASAP7_75t_R register___U13973 ( .A(register__n9340), .Y(register__n9339) );
  BUFx4f_ASAP7_75t_R register___U13974 ( .A(register__n6866), .Y(register__n9340) );
  BUFx6f_ASAP7_75t_R register___U13975 ( .A(register__n9342), .Y(register__n9341) );
  BUFx4f_ASAP7_75t_R register___U13976 ( .A(register__n8439), .Y(register__n9342) );
  BUFx6f_ASAP7_75t_R register___U13977 ( .A(register__n9344), .Y(register__n9343) );
  BUFx4f_ASAP7_75t_R register___U13978 ( .A(register__n6099), .Y(register__n9344) );
  BUFx4f_ASAP7_75t_R register___U13979 ( .A(register__n6883), .Y(register__n9346) );
  BUFx6f_ASAP7_75t_R register___U13980 ( .A(register__n9348), .Y(register__n9347) );
  BUFx4f_ASAP7_75t_R register___U13981 ( .A(register__n6886), .Y(register__n9348) );
  BUFx4f_ASAP7_75t_R register___U13982 ( .A(register__net119330), .Y(register__net93468) );
  BUFx4f_ASAP7_75t_R register___U13983 ( .A(register__net110122), .Y(register__net93464) );
  BUFx6f_ASAP7_75t_R register___U13984 ( .A(register__n9350), .Y(register__n9349) );
  BUFx4f_ASAP7_75t_R register___U13985 ( .A(register__n6935), .Y(register__n9350) );
  BUFx4f_ASAP7_75t_R register___U13986 ( .A(register__net112281), .Y(register__net93456) );
  BUFx6f_ASAP7_75t_R register___U13987 ( .A(register__n9352), .Y(register__n9351) );
  BUFx4f_ASAP7_75t_R register___U13988 ( .A(register__n7829), .Y(register__n9352) );
  BUFx6f_ASAP7_75t_R register___U13989 ( .A(register__n9354), .Y(register__n9353) );
  BUFx4f_ASAP7_75t_R register___U13990 ( .A(register__n6671), .Y(register__n9354) );
  BUFx6f_ASAP7_75t_R register___U13991 ( .A(register__n9356), .Y(register__n9355) );
  BUFx4f_ASAP7_75t_R register___U13992 ( .A(register__n6311), .Y(register__n9356) );
  BUFx4f_ASAP7_75t_R register___U13993 ( .A(register__net112533), .Y(register__net93440) );
  BUFx6f_ASAP7_75t_R register___U13994 ( .A(register__n9358), .Y(register__n9357) );
  BUFx4f_ASAP7_75t_R register___U13995 ( .A(register__n6319), .Y(register__n9358) );
  BUFx6f_ASAP7_75t_R register___U13996 ( .A(register__n9360), .Y(register__n9359) );
  BUFx4f_ASAP7_75t_R register___U13997 ( .A(register__n6084), .Y(register__n9360) );
  BUFx6f_ASAP7_75t_R register___U13998 ( .A(register__n9362), .Y(register__n9361) );
  BUFx4f_ASAP7_75t_R register___U13999 ( .A(register__n7418), .Y(register__n9362) );
  BUFx6f_ASAP7_75t_R register___U14000 ( .A(register__n9364), .Y(register__n9363) );
  BUFx4f_ASAP7_75t_R register___U14001 ( .A(register__n5865), .Y(register__n9364) );
  BUFx4f_ASAP7_75t_R register___U14002 ( .A(register__net108027), .Y(register__net93420) );
  BUFx4f_ASAP7_75t_R register___U14003 ( .A(register__n8128), .Y(register__n9366) );
  BUFx6f_ASAP7_75t_R register___U14004 ( .A(register__n9368), .Y(register__n9367) );
  BUFx4f_ASAP7_75t_R register___U14005 ( .A(register__n7802), .Y(register__n9368) );
  BUFx4f_ASAP7_75t_R register___U14006 ( .A(register__net112313), .Y(register__net93408) );
  BUFx4f_ASAP7_75t_R register___U14007 ( .A(register__net115984), .Y(register__net93404) );
  BUFx6f_ASAP7_75t_R register___U14008 ( .A(register__n9370), .Y(register__n9369) );
  BUFx4f_ASAP7_75t_R register___U14009 ( .A(register__n7198), .Y(register__n9370) );
  BUFx4f_ASAP7_75t_R register___U14010 ( .A(register__net107940), .Y(register__net93396) );
  BUFx6f_ASAP7_75t_R register___U14011 ( .A(register__n9372), .Y(register__n9371) );
  BUFx4f_ASAP7_75t_R register___U14012 ( .A(register__n6675), .Y(register__n9372) );
  BUFx6f_ASAP7_75t_R register___U14013 ( .A(register__n9374), .Y(register__n9373) );
  BUFx4f_ASAP7_75t_R register___U14014 ( .A(register__n8054), .Y(register__n9374) );
  BUFx6f_ASAP7_75t_R register___U14015 ( .A(register__n9376), .Y(register__n9375) );
  BUFx4f_ASAP7_75t_R register___U14016 ( .A(register__n8056), .Y(register__n9376) );
  BUFx6f_ASAP7_75t_R register___U14017 ( .A(register__n9378), .Y(register__n9377) );
  BUFx4f_ASAP7_75t_R register___U14018 ( .A(register__n7844), .Y(register__n9378) );
  BUFx6f_ASAP7_75t_R register___U14019 ( .A(register__net93376), .Y(register__net93375) );
  BUFx4f_ASAP7_75t_R register___U14020 ( .A(register__net103385), .Y(register__net93376) );
  INVx2_ASAP7_75t_R register___U14021 ( .A(register__n11865), .Y(register__n11863) );
  BUFx12f_ASAP7_75t_R register___U14022 ( .A(register__n3936), .Y(register__n11865) );
  BUFx6f_ASAP7_75t_R register___U14023 ( .A(register__n9381), .Y(register__n9380) );
  BUFx4f_ASAP7_75t_R register___U14024 ( .A(register__n6326), .Y(register__n9381) );
  BUFx6f_ASAP7_75t_R register___U14025 ( .A(register__n9383), .Y(register__n9382) );
  BUFx4f_ASAP7_75t_R register___U14026 ( .A(register__n6082), .Y(register__n9383) );
  BUFx6f_ASAP7_75t_R register___U14027 ( .A(register__n9385), .Y(register__n9384) );
  BUFx4f_ASAP7_75t_R register___U14028 ( .A(register__n8048), .Y(register__n9385) );
  BUFx6f_ASAP7_75t_R register___U14029 ( .A(register__n9387), .Y(register__n9386) );
  BUFx4f_ASAP7_75t_R register___U14030 ( .A(register__n6912), .Y(register__n9387) );
  BUFx6f_ASAP7_75t_R register___U14031 ( .A(register__n5347), .Y(register__n12353) );
  OA22x2_ASAP7_75t_R register___U14032 ( .A1(register__n12322), .A2(register__n4033), .B1(register__n9252), .B2(register__n11842), 
        .Y(register__n12533) );
  INVx1_ASAP7_75t_R register___U14033 ( .A(register__n6515), .Y(register__n9390) );
  OA22x2_ASAP7_75t_R register___U14034 ( .A1(register__n12080), .A2(register__n4033), .B1(register__n9341), .B2(register__n3212), 
        .Y(register__n12543) );
  INVx1_ASAP7_75t_R register___U14035 ( .A(register__n6502), .Y(register__n9391) );
  OA22x2_ASAP7_75t_R register___U14036 ( .A1(register__n12236), .A2(register__n4033), .B1(register__n9266), .B2(register__n4845), 
        .Y(register__n12536) );
  OA22x2_ASAP7_75t_R register___U14037 ( .A1(register__net64002), .A2(register__n1092), .B1(register__net93797), .B2(
        n5173), .Y(register__n13076) );
  OA22x2_ASAP7_75t_R register___U14038 ( .A1(register__n12465), .A2(register__n4033), .B1(register__n9268), .B2(register__n11920), 
        .Y(register__n12523) );
  INVx1_ASAP7_75t_R register___U14039 ( .A(register__n4525), .Y(register__n9392) );
  OA22x2_ASAP7_75t_R register___U14040 ( .A1(register__n12171), .A2(register__n4033), .B1(register__n9270), .B2(register__n5050), 
        .Y(register__n12539) );
  INVx1_ASAP7_75t_R register___U14041 ( .A(register__n4302), .Y(register__n9393) );
  OA22x2_ASAP7_75t_R register___U14042 ( .A1(register__net146308), .A2(register__n1616), .B1(register__n9274), .B2(
        n3257), .Y(register__n13069) );
  OA22x2_ASAP7_75t_R register___U14043 ( .A1(register__n12464), .A2(register__n1549), .B1(register__n9299), .B2(register__n1542), 
        .Y(register__n12580) );
  OA22x2_ASAP7_75t_R register___U14044 ( .A1(register__n12284), .A2(register__n1092), .B1(register__n9303), .B2(register__n11758), 
        .Y(register__n13073) );
  INVx1_ASAP7_75t_R register___U14045 ( .A(register__n4883), .Y(register__n9395) );
  OA22x2_ASAP7_75t_R register___U14046 ( .A1(register__net62828), .A2(register__n956), .B1(register__net96915), .B2(
        n959), .Y(register__n13011) );
  BUFx6f_ASAP7_75t_R register___U14047 ( .A(register__n12449), .Y(register__n12437) );
  BUFx6f_ASAP7_75t_R register___U14048 ( .A(register__n6269), .Y(register__n12443) );
  OA22x2_ASAP7_75t_R register___U14049 ( .A1(register__register__n11997), .A2(register__n119), .B1(register__n9256), .B2(register__n1534), 
        .Y(register__n12604) );
  OA22x2_ASAP7_75t_R register___U14050 ( .A1(register__n3593), .A2(register__n1069), .B1(register__n6321), .B2(register__n81), 
        .Y(register__n12829) );
  INVx1_ASAP7_75t_R register___U14051 ( .A(register__n3765), .Y(register__n9397) );
  OA22x2_ASAP7_75t_R register___U14052 ( .A1(register__n11990), .A2(register__n1416), .B1(register__n4959), .B2(register__n1417), 
        .Y(register__n13007) );
  INVx1_ASAP7_75t_R register___U14053 ( .A(register__n5962), .Y(register__n9398) );
  OA22x2_ASAP7_75t_R register___U14054 ( .A1(register__n3441), .A2(register__n895), .B1(register__n9258), .B2(register__n899), 
        .Y(register__n13061) );
  INVx1_ASAP7_75t_R register___U14055 ( .A(register__n8366), .Y(register__n9399) );
  OA22x2_ASAP7_75t_R register___U14056 ( .A1(register__net62820), .A2(register__n11868), .B1(register__net93661), .B2(
        n11746), .Y(register__n13264) );
  OA22x2_ASAP7_75t_R register___U14057 ( .A1(register__n12113), .A2(register__n577), .B1(register__n9319), .B2(register__n579), 
        .Y(register__n13226) );
  INVx1_ASAP7_75t_R register___U14058 ( .A(register__n5578), .Y(register__n9400) );
  OA22x2_ASAP7_75t_R register___U14059 ( .A1(register__n12404), .A2(register__n578), .B1(register__n9365), .B2(register__n586), 
        .Y(register__n13213) );
  OA22x2_ASAP7_75t_R register___U14060 ( .A1(register__net62822), .A2(register__n575), .B1(register__net93408), .B2(
        n582), .Y(register__n13210) );
  INVx1_ASAP7_75t_R register___U14061 ( .A(register__n5580), .Y(register__n9402) );
  BUFx6f_ASAP7_75t_R register___U14062 ( .A(register__net92027), .Y(register__net63270) );
  BUFx6f_ASAP7_75t_R register___U14063 ( .A(register__net92027), .Y(register__net63278) );
  OA22x2_ASAP7_75t_R register___U14064 ( .A1(register__n12256), .A2(register__n462), .B1(register__n9380), .B2(register__n465), 
        .Y(register__n12931) );
  OA22x2_ASAP7_75t_R register___U14065 ( .A1(register__n12254), .A2(register__n894), .B1(register__n9384), .B2(register__n902), 
        .Y(register__n13048) );
  BUFx12f_ASAP7_75t_R register___U14066 ( .A(register__n2963), .Y(register__n9406) );
  BUFx16f_ASAP7_75t_R register___U14067 ( .A(register__n11965), .Y(register__n11966) );
  BUFx12f_ASAP7_75t_R register___U14068 ( .A(register__net127722), .Y(register__net91940) );
  BUFx12f_ASAP7_75t_R register___U14069 ( .A(register__net64980), .Y(register__net91919) );
  BUFx12f_ASAP7_75t_R register___U14070 ( .A(register__net64958), .Y(register__net91920) );
  BUFx4f_ASAP7_75t_R register___U14071 ( .A(register__net91670), .Y(register__net114452) );
  BUFx3_ASAP7_75t_R register___U14072 ( .A(register__net114451), .Y(register__net91670) );
  BUFx4f_ASAP7_75t_R register___U14073 ( .A(register__net95070), .Y(register__net91591) );
  BUFx6f_ASAP7_75t_R register___U14074 ( .A(register__n9418), .Y(register__n9417) );
  BUFx4f_ASAP7_75t_R register___U14075 ( .A(register__n6118), .Y(register__n9418) );
  BUFx4f_ASAP7_75t_R register___U14076 ( .A(register__net112207), .Y(register__net91583) );
  BUFx6f_ASAP7_75t_R register___U14077 ( .A(register__n9420), .Y(register__n9419) );
  BUFx4f_ASAP7_75t_R register___U14078 ( .A(register__n6313), .Y(register__n9420) );
  BUFx6f_ASAP7_75t_R register___U14079 ( .A(register__n9422), .Y(register__n9421) );
  BUFx4f_ASAP7_75t_R register___U14080 ( .A(register__n7163), .Y(register__n9422) );
  BUFx6f_ASAP7_75t_R register___U14081 ( .A(register__n9426), .Y(register__n9425) );
  BUFx4f_ASAP7_75t_R register___U14082 ( .A(register__n6571), .Y(register__n9426) );
  BUFx6f_ASAP7_75t_R register___U14083 ( .A(register__n9428), .Y(register__n9427) );
  BUFx4f_ASAP7_75t_R register___U14084 ( .A(register__n6593), .Y(register__n9428) );
  BUFx6f_ASAP7_75t_R register___U14085 ( .A(register__n9430), .Y(register__n9429) );
  BUFx4f_ASAP7_75t_R register___U14086 ( .A(register__n8435), .Y(register__n9430) );
  BUFx6f_ASAP7_75t_R register___U14087 ( .A(register__n9432), .Y(register__n9431) );
  BUFx4f_ASAP7_75t_R register___U14088 ( .A(register__n8437), .Y(register__n9432) );
  BUFx6f_ASAP7_75t_R register___U14089 ( .A(register__n9436), .Y(register__n9435) );
  BUFx4f_ASAP7_75t_R register___U14090 ( .A(register__n8388), .Y(register__n9436) );
  BUFx6f_ASAP7_75t_R register___U14091 ( .A(register__n9438), .Y(register__n9437) );
  BUFx4f_ASAP7_75t_R register___U14092 ( .A(register__n8845), .Y(register__n9438) );
  BUFx6f_ASAP7_75t_R register___U14093 ( .A(register__n9440), .Y(register__n9439) );
  BUFx4f_ASAP7_75t_R register___U14094 ( .A(register__n8847), .Y(register__n9440) );
  BUFx6f_ASAP7_75t_R register___U14095 ( .A(register__net91528), .Y(register__net91527) );
  BUFx4f_ASAP7_75t_R register___U14096 ( .A(register__net98677), .Y(register__net91528) );
  BUFx4f_ASAP7_75t_R register___U14097 ( .A(register__net98673), .Y(register__net91523) );
  BUFx6f_ASAP7_75t_R register___U14098 ( .A(register__n9442), .Y(register__n9441) );
  BUFx4f_ASAP7_75t_R register___U14099 ( .A(register__n8849), .Y(register__n9442) );
  BUFx6f_ASAP7_75t_R register___U14100 ( .A(register__n9444), .Y(register__n9443) );
  BUFx4f_ASAP7_75t_R register___U14101 ( .A(register__n8390), .Y(register__n9444) );
  BUFx6f_ASAP7_75t_R register___U14102 ( .A(register__n9446), .Y(register__n9445) );
  BUFx4f_ASAP7_75t_R register___U14103 ( .A(register__n8392), .Y(register__n9446) );
  BUFx6f_ASAP7_75t_R register___U14104 ( .A(register__n9448), .Y(register__n9447) );
  BUFx4f_ASAP7_75t_R register___U14105 ( .A(register__n8851), .Y(register__n9448) );
  BUFx6f_ASAP7_75t_R register___U14106 ( .A(register__n9450), .Y(register__n9449) );
  BUFx4f_ASAP7_75t_R register___U14107 ( .A(register__n8394), .Y(register__n9450) );
  BUFx6f_ASAP7_75t_R register___U14108 ( .A(register__n9452), .Y(register__n9451) );
  BUFx4f_ASAP7_75t_R register___U14109 ( .A(register__n8853), .Y(register__n9452) );
  BUFx6f_ASAP7_75t_R register___U14110 ( .A(register__net91496), .Y(register__net91495) );
  BUFx4f_ASAP7_75t_R register___U14111 ( .A(register__net98657), .Y(register__net91496) );
  BUFx6f_ASAP7_75t_R register___U14112 ( .A(register__n9454), .Y(register__n9453) );
  BUFx4f_ASAP7_75t_R register___U14113 ( .A(register__n8855), .Y(register__n9454) );
  BUFx6f_ASAP7_75t_R register___U14114 ( .A(register__n9456), .Y(register__n9455) );
  BUFx4f_ASAP7_75t_R register___U14115 ( .A(register__n8396), .Y(register__n9456) );
  BUFx6f_ASAP7_75t_R register___U14116 ( .A(register__n9458), .Y(register__n9457) );
  BUFx4f_ASAP7_75t_R register___U14117 ( .A(register__n8398), .Y(register__n9458) );
  BUFx6f_ASAP7_75t_R register___U14118 ( .A(register__n9460), .Y(register__n9459) );
  BUFx4f_ASAP7_75t_R register___U14119 ( .A(register__n8044), .Y(register__n9460) );
  BUFx6f_ASAP7_75t_R register___U14120 ( .A(register__n9462), .Y(register__n9461) );
  BUFx4f_ASAP7_75t_R register___U14121 ( .A(register__n8402), .Y(register__n9462) );
  BUFx6f_ASAP7_75t_R register___U14122 ( .A(register__n9464), .Y(register__n9463) );
  BUFx4f_ASAP7_75t_R register___U14123 ( .A(register__n8863), .Y(register__n9464) );
  BUFx6f_ASAP7_75t_R register___U14124 ( .A(register__n9466), .Y(register__n9465) );
  BUFx4f_ASAP7_75t_R register___U14125 ( .A(register__n8865), .Y(register__n9466) );
  BUFx4f_ASAP7_75t_R register___U14126 ( .A(register__net98637), .Y(register__net91463) );
  BUFx6f_ASAP7_75t_R register___U14127 ( .A(register__n9468), .Y(register__n9467) );
  BUFx4f_ASAP7_75t_R register___U14128 ( .A(register__n8867), .Y(register__n9468) );
  BUFx6f_ASAP7_75t_R register___U14129 ( .A(register__n9470), .Y(register__n9469) );
  BUFx4f_ASAP7_75t_R register___U14130 ( .A(register__n8046), .Y(register__n9470) );
  BUFx6f_ASAP7_75t_R register___U14131 ( .A(register__n9472), .Y(register__n9471) );
  BUFx4f_ASAP7_75t_R register___U14132 ( .A(register__n8881), .Y(register__n9472) );
  BUFx6f_ASAP7_75t_R register___U14133 ( .A(register__net91448), .Y(register__net91447) );
  BUFx4f_ASAP7_75t_R register___U14134 ( .A(register__net101305), .Y(register__net91448) );
  BUFx6f_ASAP7_75t_R register___U14135 ( .A(register__n9474), .Y(register__n9473) );
  BUFx4f_ASAP7_75t_R register___U14136 ( .A(register__n7745), .Y(register__n9474) );
  BUFx6f_ASAP7_75t_R register___U14137 ( .A(register__n9476), .Y(register__n9475) );
  BUFx4f_ASAP7_75t_R register___U14138 ( .A(register__n8058), .Y(register__n9476) );
  BUFx6f_ASAP7_75t_R register___U14139 ( .A(register__n9478), .Y(register__n9477) );
  BUFx4f_ASAP7_75t_R register___U14140 ( .A(register__n7761), .Y(register__n9478) );
  BUFx6f_ASAP7_75t_R register___U14141 ( .A(register__n9480), .Y(register__n9479) );
  BUFx4f_ASAP7_75t_R register___U14142 ( .A(register__n8410), .Y(register__n9480) );
  BUFx6f_ASAP7_75t_R register___U14143 ( .A(register__n9482), .Y(register__n9481) );
  BUFx4f_ASAP7_75t_R register___U14144 ( .A(register__n8887), .Y(register__n9482) );
  BUFx6f_ASAP7_75t_R register___U14145 ( .A(register__n9484), .Y(register__n9483) );
  BUFx4f_ASAP7_75t_R register___U14146 ( .A(register__n8060), .Y(register__n9484) );
  BUFx6f_ASAP7_75t_R register___U14147 ( .A(register__n9486), .Y(register__n9485) );
  BUFx4f_ASAP7_75t_R register___U14148 ( .A(register__n8412), .Y(register__n9486) );
  BUFx6f_ASAP7_75t_R register___U14149 ( .A(register__n9488), .Y(register__n9487) );
  BUFx4f_ASAP7_75t_R register___U14150 ( .A(register__n8417), .Y(register__n9488) );
  BUFx6f_ASAP7_75t_R register___U14151 ( .A(register__n9490), .Y(register__n9489) );
  BUFx4f_ASAP7_75t_R register___U14152 ( .A(register__n8419), .Y(register__n9490) );
  BUFx6f_ASAP7_75t_R register___U14153 ( .A(register__n9492), .Y(register__n9491) );
  BUFx4f_ASAP7_75t_R register___U14154 ( .A(register__n8902), .Y(register__n9492) );
  BUFx6f_ASAP7_75t_R register___U14155 ( .A(register__n9494), .Y(register__n9493) );
  BUFx4f_ASAP7_75t_R register___U14156 ( .A(register__n8421), .Y(register__n9494) );
  BUFx6f_ASAP7_75t_R register___U14157 ( .A(register__n9496), .Y(register__n9495) );
  BUFx4f_ASAP7_75t_R register___U14158 ( .A(register__n8904), .Y(register__n9496) );
  BUFx6f_ASAP7_75t_R register___U14159 ( .A(register__net91396), .Y(register__net91395) );
  BUFx4f_ASAP7_75t_R register___U14160 ( .A(register__net98582), .Y(register__net91396) );
  BUFx6f_ASAP7_75t_R register___U14161 ( .A(register__n9498), .Y(register__n9497) );
  BUFx4f_ASAP7_75t_R register___U14162 ( .A(register__n8906), .Y(register__n9498) );
  BUFx6f_ASAP7_75t_R register___U14163 ( .A(register__n9500), .Y(register__n9499) );
  BUFx4f_ASAP7_75t_R register___U14164 ( .A(register__n8423), .Y(register__n9500) );
  BUFx6f_ASAP7_75t_R register___U14165 ( .A(register__n9502), .Y(register__n9501) );
  BUFx4f_ASAP7_75t_R register___U14166 ( .A(register__n8425), .Y(register__n9502) );
  BUFx6f_ASAP7_75t_R register___U14167 ( .A(register__n9504), .Y(register__n9503) );
  BUFx4f_ASAP7_75t_R register___U14168 ( .A(register__n8433), .Y(register__n9504) );
  BUFx6f_ASAP7_75t_R register___U14169 ( .A(register__net91376), .Y(register__net91375) );
  BUFx4f_ASAP7_75t_R register___U14170 ( .A(register__net98530), .Y(register__net91376) );
  BUFx6f_ASAP7_75t_R register___U14171 ( .A(register__n9506), .Y(register__n9505) );
  BUFx4f_ASAP7_75t_R register___U14172 ( .A(register__n8964), .Y(register__n9506) );
  BUFx6f_ASAP7_75t_R register___U14173 ( .A(register__net91368), .Y(register__net91367) );
  BUFx4f_ASAP7_75t_R register___U14174 ( .A(register__net98526), .Y(register__net91368) );
  BUFx6f_ASAP7_75t_R register___U14175 ( .A(register__n9508), .Y(register__n9507) );
  BUFx4f_ASAP7_75t_R register___U14176 ( .A(register__n8969), .Y(register__n9508) );
  BUFx6f_ASAP7_75t_R register___U14177 ( .A(register__n9510), .Y(register__n9509) );
  BUFx4f_ASAP7_75t_R register___U14178 ( .A(register__n8974), .Y(register__n9510) );
  BUFx6f_ASAP7_75t_R register___U14179 ( .A(register__n9512), .Y(register__n9511) );
  BUFx4f_ASAP7_75t_R register___U14180 ( .A(register__n8976), .Y(register__n9512) );
  BUFx6f_ASAP7_75t_R register___U14181 ( .A(register__net91348), .Y(register__net91347) );
  BUFx4f_ASAP7_75t_R register___U14182 ( .A(register__net103622), .Y(register__net91348) );
  BUFx6f_ASAP7_75t_R register___U14183 ( .A(register__n9516), .Y(register__n9515) );
  BUFx4f_ASAP7_75t_R register___U14184 ( .A(register__n8984), .Y(register__n9516) );
  BUFx4f_ASAP7_75t_R register___U14185 ( .A(register__net98518), .Y(register__net91335) );
  BUFx6f_ASAP7_75t_R register___U14186 ( .A(register__n9520), .Y(register__n9519) );
  BUFx4f_ASAP7_75t_R register___U14187 ( .A(register__n8993), .Y(register__n9520) );
  BUFx6f_ASAP7_75t_R register___U14188 ( .A(register__n9526), .Y(register__n9525) );
  BUFx4f_ASAP7_75t_R register___U14189 ( .A(register__n8100), .Y(register__n9526) );
  BUFx4f_ASAP7_75t_R register___U14190 ( .A(register__n7777), .Y(register__n9528) );
  BUFx6f_ASAP7_75t_R register___U14191 ( .A(register__net91308), .Y(register__net91307) );
  BUFx4f_ASAP7_75t_R register___U14192 ( .A(register__net95194), .Y(register__net91308) );
  BUFx6f_ASAP7_75t_R register___U14193 ( .A(register__n9530), .Y(register__n9529) );
  BUFx4f_ASAP7_75t_R register___U14194 ( .A(register__n8441), .Y(register__n9530) );
  BUFx6f_ASAP7_75t_R register___U14195 ( .A(register__n9532), .Y(register__n9531) );
  BUFx4f_ASAP7_75t_R register___U14196 ( .A(register__n7781), .Y(register__n9532) );
  BUFx6f_ASAP7_75t_R register___U14197 ( .A(register__n9534), .Y(register__n9533) );
  BUFx4f_ASAP7_75t_R register___U14198 ( .A(register__n9010), .Y(register__n9534) );
  BUFx6f_ASAP7_75t_R register___U14199 ( .A(register__n9536), .Y(register__n9535) );
  BUFx4f_ASAP7_75t_R register___U14200 ( .A(register__n8443), .Y(register__n9536) );
  BUFx6f_ASAP7_75t_R register___U14201 ( .A(register__n9538), .Y(register__n9537) );
  BUFx4f_ASAP7_75t_R register___U14202 ( .A(register__n9012), .Y(register__n9538) );
  BUFx6f_ASAP7_75t_R register___U14203 ( .A(register__n9540), .Y(register__n9539) );
  BUFx4f_ASAP7_75t_R register___U14204 ( .A(register__n8448), .Y(register__n9540) );
  BUFx6f_ASAP7_75t_R register___U14205 ( .A(register__n9542), .Y(register__n9541) );
  BUFx4f_ASAP7_75t_R register___U14206 ( .A(register__n8450), .Y(register__n9542) );
  BUFx6f_ASAP7_75t_R register___U14207 ( .A(register__n9544), .Y(register__n9543) );
  BUFx4f_ASAP7_75t_R register___U14208 ( .A(register__n9022), .Y(register__n9544) );
  BUFx6f_ASAP7_75t_R register___U14209 ( .A(register__n9546), .Y(register__n9545) );
  BUFx4f_ASAP7_75t_R register___U14210 ( .A(register__n9029), .Y(register__n9546) );
  BUFx6f_ASAP7_75t_R register___U14211 ( .A(register__n9548), .Y(register__n9547) );
  BUFx4f_ASAP7_75t_R register___U14212 ( .A(register__n9031), .Y(register__n9548) );
  BUFx6f_ASAP7_75t_R register___U14213 ( .A(register__net91264), .Y(register__net91263) );
  BUFx4f_ASAP7_75t_R register___U14214 ( .A(register__net103580), .Y(register__net91264) );
  BUFx4f_ASAP7_75t_R register___U14215 ( .A(register__net95118), .Y(register__net91259) );
  BUFx4f_ASAP7_75t_R register___U14216 ( .A(register__net95114), .Y(register__net91255) );
  BUFx6f_ASAP7_75t_R register___U14217 ( .A(register__n9550), .Y(register__n9549) );
  BUFx4f_ASAP7_75t_R register___U14218 ( .A(register__n8459), .Y(register__n9550) );
  BUFx6f_ASAP7_75t_R register___U14219 ( .A(register__n9552), .Y(register__n9551) );
  BUFx4f_ASAP7_75t_R register___U14220 ( .A(register__n9039), .Y(register__n9552) );
  BUFx6f_ASAP7_75t_R register___U14221 ( .A(register__n9554), .Y(register__n9553) );
  BUFx4f_ASAP7_75t_R register___U14222 ( .A(register__n8463), .Y(register__n9554) );
  BUFx6f_ASAP7_75t_R register___U14223 ( .A(register__n9556), .Y(register__n9555) );
  BUFx4f_ASAP7_75t_R register___U14224 ( .A(register__n8465), .Y(register__n9556) );
  BUFx6f_ASAP7_75t_R register___U14225 ( .A(register__n9558), .Y(register__n9557) );
  BUFx4f_ASAP7_75t_R register___U14226 ( .A(register__n8467), .Y(register__n9558) );
  BUFx6f_ASAP7_75t_R register___U14227 ( .A(register__n9560), .Y(register__n9559) );
  BUFx4f_ASAP7_75t_R register___U14228 ( .A(register__n8469), .Y(register__n9560) );
  BUFx6f_ASAP7_75t_R register___U14229 ( .A(register__n9562), .Y(register__n9561) );
  BUFx4f_ASAP7_75t_R register___U14230 ( .A(register__n7790), .Y(register__n9562) );
  BUFx6f_ASAP7_75t_R register___U14231 ( .A(register__n9564), .Y(register__n9563) );
  BUFx4f_ASAP7_75t_R register___U14232 ( .A(register__n7792), .Y(register__n9564) );
  BUFx4f_ASAP7_75t_R register___U14233 ( .A(register__net103540), .Y(register__net91220) );
  BUFx6f_ASAP7_75t_R register___U14234 ( .A(register__n9566), .Y(register__n9565) );
  BUFx4f_ASAP7_75t_R register___U14235 ( .A(register__n9046), .Y(register__n9566) );
  BUFx6f_ASAP7_75t_R register___U14236 ( .A(register__n9568), .Y(register__n9567) );
  BUFx4f_ASAP7_75t_R register___U14237 ( .A(register__n7796), .Y(register__n9568) );
  BUFx6f_ASAP7_75t_R register___U14238 ( .A(register__n9570), .Y(register__n9569) );
  BUFx4f_ASAP7_75t_R register___U14239 ( .A(register__n7804), .Y(register__n9570) );
  BUFx6f_ASAP7_75t_R register___U14240 ( .A(register__net91204), .Y(register__net91203) );
  BUFx4f_ASAP7_75t_R register___U14241 ( .A(register__net95048), .Y(register__net91204) );
  BUFx6f_ASAP7_75t_R register___U14242 ( .A(register__n9572), .Y(register__n9571) );
  BUFx4f_ASAP7_75t_R register___U14243 ( .A(register__n8149), .Y(register__n9572) );
  BUFx6f_ASAP7_75t_R register___U14244 ( .A(register__n9574), .Y(register__n9573) );
  BUFx4f_ASAP7_75t_R register___U14245 ( .A(register__n6833), .Y(register__n9574) );
  BUFx4f_ASAP7_75t_R register___U14246 ( .A(register__net103751), .Y(register__net91105) );
  BUFx6f_ASAP7_75t_R register___U14247 ( .A(register__n9576), .Y(register__n9575) );
  BUFx4f_ASAP7_75t_R register___U14248 ( .A(register__n6060), .Y(register__n9576) );
  BUFx6f_ASAP7_75t_R register___U14249 ( .A(register__n9578), .Y(register__n9577) );
  BUFx4f_ASAP7_75t_R register___U14250 ( .A(register__n6062), .Y(register__n9578) );
  BUFx6f_ASAP7_75t_R register___U14251 ( .A(register__n9580), .Y(register__n9579) );
  BUFx4f_ASAP7_75t_R register___U14252 ( .A(register__n5186), .Y(register__n9580) );
  BUFx6f_ASAP7_75t_R register___U14253 ( .A(register__n9582), .Y(register__n9581) );
  BUFx4f_ASAP7_75t_R register___U14254 ( .A(register__n7397), .Y(register__n9582) );
  BUFx6f_ASAP7_75t_R register___U14255 ( .A(register__n9584), .Y(register__n9583) );
  BUFx4f_ASAP7_75t_R register___U14256 ( .A(register__n5188), .Y(register__n9584) );
  BUFx6f_ASAP7_75t_R register___U14257 ( .A(register__n9586), .Y(register__n9585) );
  BUFx4f_ASAP7_75t_R register___U14258 ( .A(register__n5193), .Y(register__n9586) );
  BUFx4f_ASAP7_75t_R register___U14259 ( .A(register__n7729), .Y(register__n9588) );
  BUFx4f_ASAP7_75t_R register___U14260 ( .A(register__net101357), .Y(register__net91073) );
  BUFx4f_ASAP7_75t_R register___U14261 ( .A(register__net123675), .Y(register__net91069) );
  BUFx6f_ASAP7_75t_R register___U14262 ( .A(register__n9590), .Y(register__n9589) );
  BUFx4f_ASAP7_75t_R register___U14263 ( .A(register__n6064), .Y(register__n9590) );
  BUFx6f_ASAP7_75t_R register___U14264 ( .A(register__n9592), .Y(register__n9591) );
  BUFx4f_ASAP7_75t_R register___U14265 ( .A(register__n8384), .Y(register__n9592) );
  BUFx6f_ASAP7_75t_R register___U14266 ( .A(register__n9594), .Y(register__n9593) );
  BUFx4f_ASAP7_75t_R register___U14267 ( .A(register__n7402), .Y(register__n9594) );
  BUFx6f_ASAP7_75t_R register___U14268 ( .A(register__n9596), .Y(register__n9595) );
  BUFx4f_ASAP7_75t_R register___U14269 ( .A(register__n6066), .Y(register__n9596) );
  BUFx6f_ASAP7_75t_R register___U14270 ( .A(register__n9598), .Y(register__n9597) );
  BUFx4f_ASAP7_75t_R register___U14271 ( .A(register__n5361), .Y(register__n9598) );
  BUFx6f_ASAP7_75t_R register___U14272 ( .A(register__net91046), .Y(register__net91045) );
  BUFx4f_ASAP7_75t_R register___U14273 ( .A(register__net98689), .Y(register__net91046) );
  BUFx6f_ASAP7_75t_R register___U14274 ( .A(register__n9600), .Y(register__n9599) );
  BUFx4f_ASAP7_75t_R register___U14275 ( .A(register__n7406), .Y(register__n9600) );
  BUFx6f_ASAP7_75t_R register___U14276 ( .A(register__n9602), .Y(register__n9601) );
  BUFx4f_ASAP7_75t_R register___U14277 ( .A(register__n6068), .Y(register__n9602) );
  BUFx4f_ASAP7_75t_R register___U14278 ( .A(register__net108118), .Y(register__net91033) );
  BUFx6f_ASAP7_75t_R register___U14279 ( .A(register__n9604), .Y(register__n9603) );
  BUFx4f_ASAP7_75t_R register___U14280 ( .A(register__n7732), .Y(register__n9604) );
  BUFx6f_ASAP7_75t_R register___U14281 ( .A(register__n9606), .Y(register__n9605) );
  BUFx4f_ASAP7_75t_R register___U14282 ( .A(register__n8386), .Y(register__n9606) );
  BUFx6f_ASAP7_75t_R register___U14283 ( .A(register__n9608), .Y(register__n9607) );
  BUFx4f_ASAP7_75t_R register___U14284 ( .A(register__n6835), .Y(register__n9608) );
  BUFx6f_ASAP7_75t_R register___U14285 ( .A(register__n9610), .Y(register__n9609) );
  BUFx4f_ASAP7_75t_R register___U14286 ( .A(register__n6840), .Y(register__n9610) );
  BUFx4f_ASAP7_75t_R register___U14287 ( .A(register__net116110), .Y(register__net91001) );
  BUFx4f_ASAP7_75t_R register___U14288 ( .A(register__net112549), .Y(register__net90997) );
  BUFx6f_ASAP7_75t_R register___U14289 ( .A(register__n9616), .Y(register__n9615) );
  BUFx4f_ASAP7_75t_R register___U14290 ( .A(register__n6074), .Y(register__n9616) );
  BUFx6f_ASAP7_75t_R register___U14291 ( .A(register__n9618), .Y(register__n9617) );
  BUFx4f_ASAP7_75t_R register___U14292 ( .A(register__n6076), .Y(register__n9618) );
  BUFx6f_ASAP7_75t_R register___U14293 ( .A(register__n9620), .Y(register__n9619) );
  BUFx4f_ASAP7_75t_R register___U14294 ( .A(register__n6078), .Y(register__n9620) );
  BUFx6f_ASAP7_75t_R register___U14295 ( .A(register__n9622), .Y(register__n9621) );
  BUFx4f_ASAP7_75t_R register___U14296 ( .A(register__n6305), .Y(register__n9622) );
  BUFx6f_ASAP7_75t_R register___U14297 ( .A(register__n9624), .Y(register__n9623) );
  BUFx4f_ASAP7_75t_R register___U14298 ( .A(register__n5669), .Y(register__n9624) );
  BUFx6f_ASAP7_75t_R register___U14299 ( .A(register__n9626), .Y(register__n9625) );
  BUFx4f_ASAP7_75t_R register___U14300 ( .A(register__n5857), .Y(register__n9626) );
  BUFx4f_ASAP7_75t_R register___U14301 ( .A(register__net117775), .Y(register__net90965) );
  BUFx4f_ASAP7_75t_R register___U14302 ( .A(register__net112541), .Y(register__net90961) );
  BUFx6f_ASAP7_75t_R register___U14303 ( .A(register__n9629), .Y(register__n9628) );
  BUFx4f_ASAP7_75t_R register___U14304 ( .A(register__n6552), .Y(register__n9629) );
  BUFx6f_ASAP7_75t_R register___U14305 ( .A(register__n9631), .Y(register__n9630) );
  BUFx4f_ASAP7_75t_R register___U14306 ( .A(register__n6844), .Y(register__n9631) );
  BUFx6f_ASAP7_75t_R register___U14307 ( .A(register__n9633), .Y(register__n9632) );
  BUFx4f_ASAP7_75t_R register___U14308 ( .A(register__n6307), .Y(register__n9633) );
  BUFx6f_ASAP7_75t_R register___U14309 ( .A(register__n9635), .Y(register__n9634) );
  BUFx4f_ASAP7_75t_R register___U14310 ( .A(register__n6309), .Y(register__n9635) );
  BUFx6f_ASAP7_75t_R register___U14311 ( .A(register__n9637), .Y(register__n9636) );
  BUFx4f_ASAP7_75t_R register___U14312 ( .A(register__n7439), .Y(register__n9637) );
  BUFx4f_ASAP7_75t_R register___U14313 ( .A(register__net116074), .Y(register__net90937) );
  BUFx6f_ASAP7_75t_R register___U14314 ( .A(register__n9639), .Y(register__n9638) );
  BUFx4f_ASAP7_75t_R register___U14315 ( .A(register__n7165), .Y(register__n9639) );
  BUFx6f_ASAP7_75t_R register___U14316 ( .A(register__n9641), .Y(register__n9640) );
  BUFx4f_ASAP7_75t_R register___U14317 ( .A(register__n8869), .Y(register__n9641) );
  BUFx4f_ASAP7_75t_R register___U14318 ( .A(register__net95618), .Y(register__net90925) );
  BUFx6f_ASAP7_75t_R register___U14319 ( .A(register__n9643), .Y(register__n9642) );
  BUFx4f_ASAP7_75t_R register___U14320 ( .A(register__n8871), .Y(register__n9643) );
  BUFx6f_ASAP7_75t_R register___U14321 ( .A(register__n9645), .Y(register__n9644) );
  BUFx4f_ASAP7_75t_R register___U14322 ( .A(register__n6573), .Y(register__n9645) );
  BUFx6f_ASAP7_75t_R register___U14323 ( .A(register__n9647), .Y(register__n9646) );
  BUFx4f_ASAP7_75t_R register___U14324 ( .A(register__n6575), .Y(register__n9647) );
  BUFx6f_ASAP7_75t_R register___U14325 ( .A(register__n9649), .Y(register__n9648) );
  BUFx4f_ASAP7_75t_R register___U14326 ( .A(register__n6336), .Y(register__n9649) );
  BUFx4f_ASAP7_75t_R register___U14327 ( .A(register__net114228), .Y(register__net90905) );
  BUFx4f_ASAP7_75t_R register___U14328 ( .A(register__net114224), .Y(register__net90901) );
  BUFx6f_ASAP7_75t_R register___U14329 ( .A(register__n9651), .Y(register__n9650) );
  BUFx4f_ASAP7_75t_R register___U14330 ( .A(register__n4378), .Y(register__n9651) );
  BUFx6f_ASAP7_75t_R register___U14331 ( .A(register__n9653), .Y(register__n9652) );
  BUFx4f_ASAP7_75t_R register___U14332 ( .A(register__n6338), .Y(register__n9653) );
  BUFx6f_ASAP7_75t_R register___U14333 ( .A(register__n9655), .Y(register__n9654) );
  BUFx4f_ASAP7_75t_R register___U14334 ( .A(register__n7167), .Y(register__n9655) );
  BUFx6f_ASAP7_75t_R register___U14335 ( .A(register__n9657), .Y(register__n9656) );
  BUFx4f_ASAP7_75t_R register___U14336 ( .A(register__n7169), .Y(register__n9657) );
  BUFx6f_ASAP7_75t_R register___U14337 ( .A(register__n9659), .Y(register__n9658) );
  BUFx4f_ASAP7_75t_R register___U14338 ( .A(register__n7171), .Y(register__n9659) );
  BUFx4f_ASAP7_75t_R register___U14339 ( .A(register__net98633), .Y(register__net90877) );
  BUFx6f_ASAP7_75t_R register___U14340 ( .A(register__n9661), .Y(register__n9660) );
  BUFx4f_ASAP7_75t_R register___U14341 ( .A(register__n7173), .Y(register__n9661) );
  BUFx6f_ASAP7_75t_R register___U14342 ( .A(register__n9663), .Y(register__n9662) );
  BUFx4f_ASAP7_75t_R register___U14343 ( .A(register__n8404), .Y(register__n9663) );
  BUFx4f_ASAP7_75t_R register___U14344 ( .A(register__net103720), .Y(register__net90865) );
  BUFx6f_ASAP7_75t_R register___U14345 ( .A(register__n9665), .Y(register__n9664) );
  BUFx4f_ASAP7_75t_R register___U14346 ( .A(register__n7741), .Y(register__n9665) );
  BUFx6f_ASAP7_75t_R register___U14347 ( .A(register__n9667), .Y(register__n9666) );
  BUFx4f_ASAP7_75t_R register___U14348 ( .A(register__n7175), .Y(register__n9667) );
  BUFx4f_ASAP7_75t_R register___U14349 ( .A(register__net101325), .Y(register__net90853) );
  BUFx6f_ASAP7_75t_R register___U14350 ( .A(register__n9669), .Y(register__n9668) );
  BUFx4f_ASAP7_75t_R register___U14351 ( .A(register__n8050), .Y(register__n9669) );
  BUFx6f_ASAP7_75t_R register___U14352 ( .A(register__n9671), .Y(register__n9670) );
  BUFx4f_ASAP7_75t_R register___U14353 ( .A(register__n8875), .Y(register__n9671) );
  BUFx6f_ASAP7_75t_R register___U14354 ( .A(register__n9673), .Y(register__n9672) );
  BUFx4f_ASAP7_75t_R register___U14355 ( .A(register__n8877), .Y(register__n9673) );
  BUFx4f_ASAP7_75t_R register___U14356 ( .A(register__n8879), .Y(register__n9675) );
  BUFx4f_ASAP7_75t_R register___U14357 ( .A(register__net101313), .Y(register__net90833) );
  BUFx4f_ASAP7_75t_R register___U14358 ( .A(register__net95594), .Y(register__net90829) );
  BUFx6f_ASAP7_75t_R register___U14359 ( .A(register__n9677), .Y(register__n9676) );
  BUFx4f_ASAP7_75t_R register___U14360 ( .A(register__n6864), .Y(register__n9677) );
  BUFx6f_ASAP7_75t_R register___U14361 ( .A(register__n9679), .Y(register__n9678) );
  BUFx4f_ASAP7_75t_R register___U14362 ( .A(register__n6577), .Y(register__n9679) );
  BUFx6f_ASAP7_75t_R register___U14363 ( .A(register__n9681), .Y(register__n9680) );
  BUFx4f_ASAP7_75t_R register___U14364 ( .A(register__n7441), .Y(register__n9681) );
  BUFx4f_ASAP7_75t_R register___U14365 ( .A(register__net98621), .Y(register__net90813) );
  BUFx6f_ASAP7_75t_R register___U14366 ( .A(register__n9683), .Y(register__n9682) );
  BUFx4f_ASAP7_75t_R register___U14367 ( .A(register__n7747), .Y(register__n9683) );
  BUFx6f_ASAP7_75t_R register___U14368 ( .A(register__n9685), .Y(register__n9684) );
  BUFx4f_ASAP7_75t_R register___U14369 ( .A(register__n7749), .Y(register__n9685) );
  BUFx6f_ASAP7_75t_R register___U14370 ( .A(register__n9687), .Y(register__n9686) );
  BUFx4f_ASAP7_75t_R register___U14371 ( .A(register__n8408), .Y(register__n9687) );
  BUFx6f_ASAP7_75t_R register___U14372 ( .A(register__n9689), .Y(register__n9688) );
  BUFx4f_ASAP7_75t_R register___U14373 ( .A(register__n7751), .Y(register__n9689) );
  BUFx4f_ASAP7_75t_R register___U14374 ( .A(register__net140427), .Y(register__net90789) );
  BUFx6f_ASAP7_75t_R register___U14375 ( .A(register__n9691), .Y(register__n9690) );
  BUFx4f_ASAP7_75t_R register___U14376 ( .A(register__n7755), .Y(register__n9691) );
  BUFx6f_ASAP7_75t_R register___U14377 ( .A(register__n9693), .Y(register__n9692) );
  BUFx4f_ASAP7_75t_R register___U14378 ( .A(register__n3691), .Y(register__n9693) );
  BUFx6f_ASAP7_75t_R register___U14379 ( .A(register__n9695), .Y(register__n9694) );
  BUFx4f_ASAP7_75t_R register___U14380 ( .A(register__n7757), .Y(register__n9695) );
  BUFx6f_ASAP7_75t_R register___U14381 ( .A(register__n9697), .Y(register__n9696) );
  BUFx4f_ASAP7_75t_R register___U14382 ( .A(register__n7759), .Y(register__n9697) );
  BUFx6f_ASAP7_75t_R register___U14383 ( .A(register__n9699), .Y(register__n9698) );
  BUFx4f_ASAP7_75t_R register___U14384 ( .A(register__n8908), .Y(register__n9699) );
  BUFx4f_ASAP7_75t_R register___U14385 ( .A(register__n8913), .Y(register__n9701) );
  BUFx4f_ASAP7_75t_R register___U14386 ( .A(register__net95498), .Y(register__net90762) );
  BUFx6f_ASAP7_75t_R register___U14387 ( .A(register__n9703), .Y(register__n9702) );
  BUFx4f_ASAP7_75t_R register___U14388 ( .A(register__n8916), .Y(register__n9703) );
  BUFx4f_ASAP7_75t_R register___U14389 ( .A(register__n8918), .Y(register__n9705) );
  BUFx4f_ASAP7_75t_R register___U14390 ( .A(register__n8924), .Y(register__n9707) );
  BUFx6f_ASAP7_75t_R register___U14391 ( .A(register__n9709), .Y(register__n9708) );
  BUFx4f_ASAP7_75t_R register___U14392 ( .A(register__n8927), .Y(register__n9709) );
  BUFx6f_ASAP7_75t_R register___U14393 ( .A(register__n9711), .Y(register__n9710) );
  BUFx4f_ASAP7_75t_R register___U14394 ( .A(register__n8932), .Y(register__n9711) );
  BUFx6f_ASAP7_75t_R register___U14395 ( .A(register__n9713), .Y(register__n9712) );
  BUFx4f_ASAP7_75t_R register___U14396 ( .A(register__n8427), .Y(register__n9713) );
  BUFx4f_ASAP7_75t_R register___U14397 ( .A(register__net95449), .Y(register__net90733) );
  BUFx4f_ASAP7_75t_R register___U14398 ( .A(register__net95442), .Y(register__net90730) );
  BUFx4f_ASAP7_75t_R register___U14399 ( .A(register__n8934), .Y(register__n9715) );
  BUFx6f_ASAP7_75t_R register___U14400 ( .A(register__n9717), .Y(register__n9716) );
  BUFx4f_ASAP7_75t_R register___U14401 ( .A(register__n7451), .Y(register__n9717) );
  BUFx6f_ASAP7_75t_R register___U14402 ( .A(register__n9719), .Y(register__n9718) );
  BUFx4f_ASAP7_75t_R register___U14403 ( .A(register__n7491), .Y(register__n9719) );
  BUFx6f_ASAP7_75t_R register___U14404 ( .A(register__n9723), .Y(register__n9722) );
  BUFx4f_ASAP7_75t_R register___U14405 ( .A(register__n6872), .Y(register__n9723) );
  BUFx4f_ASAP7_75t_R register___U14406 ( .A(register__n8971), .Y(register__n9725) );
  BUFx6f_ASAP7_75t_R register___U14407 ( .A(register__n9727), .Y(register__n9726) );
  BUFx4f_ASAP7_75t_R register___U14408 ( .A(register__n8982), .Y(register__n9727) );
  BUFx6f_ASAP7_75t_R register___U14409 ( .A(register__n9729), .Y(register__n9728) );
  BUFx4f_ASAP7_75t_R register___U14410 ( .A(register__n6350), .Y(register__n9729) );
  BUFx4f_ASAP7_75t_R register___U14411 ( .A(register__net108019), .Y(register__net90681) );
  BUFx4f_ASAP7_75t_R register___U14412 ( .A(register__net95241), .Y(register__net90677) );
  BUFx4f_ASAP7_75t_R register___U14413 ( .A(register__net105794), .Y(register__net90674) );
  BUFx4f_ASAP7_75t_R register___U14414 ( .A(register__net95234), .Y(register__net90670) );
  BUFx4f_ASAP7_75t_R register___U14415 ( .A(register__net105790), .Y(register__net90661) );
  BUFx4f_ASAP7_75t_R register___U14416 ( .A(register__net141142), .Y(register__net90657) );
  BUFx6f_ASAP7_75t_R register___U14417 ( .A(register__n9731), .Y(register__n9730) );
  BUFx4f_ASAP7_75t_R register___U14418 ( .A(register__n4969), .Y(register__n9731) );
  BUFx4f_ASAP7_75t_R register___U14419 ( .A(register__net114168), .Y(register__net90649) );
  BUFx6f_ASAP7_75t_R register___U14420 ( .A(register__n9735), .Y(register__n9734) );
  BUFx4f_ASAP7_75t_R register___U14421 ( .A(register__n6360), .Y(register__n9735) );
  BUFx4f_ASAP7_75t_R register___U14422 ( .A(register__net140415), .Y(register__net90637) );
  BUFx6f_ASAP7_75t_R register___U14423 ( .A(register__n9737), .Y(register__n9736) );
  BUFx4f_ASAP7_75t_R register___U14424 ( .A(register__n6362), .Y(register__n9737) );
  BUFx4f_ASAP7_75t_R register___U14425 ( .A(register__net116024), .Y(register__net90629) );
  BUFx6f_ASAP7_75t_R register___U14426 ( .A(register__n9741), .Y(register__n9740) );
  BUFx4f_ASAP7_75t_R register___U14427 ( .A(register__n8102), .Y(register__n9741) );
  BUFx6f_ASAP7_75t_R register___U14428 ( .A(register__n9743), .Y(register__n9742) );
  BUFx4f_ASAP7_75t_R register___U14429 ( .A(register__n5873), .Y(register__n9743) );
  BUFx6f_ASAP7_75t_R register___U14430 ( .A(register__n9747), .Y(register__n9746) );
  BUFx4f_ASAP7_75t_R register___U14431 ( .A(register__n7493), .Y(register__n9747) );
  BUFx4f_ASAP7_75t_R register___U14432 ( .A(register__n9005), .Y(register__n9749) );
  BUFx6f_ASAP7_75t_R register___U14433 ( .A(register__n9751), .Y(register__n9750) );
  BUFx4f_ASAP7_75t_R register___U14434 ( .A(register__n7185), .Y(register__n9751) );
  BUFx6f_ASAP7_75t_R register___U14435 ( .A(register__n9753), .Y(register__n9752) );
  BUFx4f_ASAP7_75t_R register___U14436 ( .A(register__n7495), .Y(register__n9753) );
  BUFx6f_ASAP7_75t_R register___U14437 ( .A(register__n9757), .Y(register__n9756) );
  BUFx4f_ASAP7_75t_R register___U14438 ( .A(register__n7785), .Y(register__n9757) );
  BUFx6f_ASAP7_75t_R register___U14439 ( .A(register__n9759), .Y(register__n9758) );
  BUFx4f_ASAP7_75t_R register___U14440 ( .A(register__n7499), .Y(register__n9759) );
  BUFx4f_ASAP7_75t_R register___U14441 ( .A(register__n7787), .Y(register__n9763) );
  BUFx6f_ASAP7_75t_R register___U14442 ( .A(register__n9765), .Y(register__n9764) );
  BUFx4f_ASAP7_75t_R register___U14443 ( .A(register__n6369), .Y(register__n9765) );
  BUFx6f_ASAP7_75t_R register___U14444 ( .A(register__n9767), .Y(register__n9766) );
  BUFx4f_ASAP7_75t_R register___U14445 ( .A(register__n7501), .Y(register__n9767) );
  BUFx6f_ASAP7_75t_R register___U14446 ( .A(register__n9769), .Y(register__n9768) );
  BUFx4f_ASAP7_75t_R register___U14447 ( .A(register__n7503), .Y(register__n9769) );
  BUFx4f_ASAP7_75t_R register___U14448 ( .A(register__n9033), .Y(register__n9771) );
  BUFx6f_ASAP7_75t_R register___U14449 ( .A(register__n9773), .Y(register__n9772) );
  BUFx4f_ASAP7_75t_R register___U14450 ( .A(register__n7189), .Y(register__n9773) );
  BUFx6f_ASAP7_75t_R register___U14451 ( .A(register__n9777), .Y(register__n9776) );
  BUFx4f_ASAP7_75t_R register___U14452 ( .A(register__n6921), .Y(register__n9777) );
  BUFx4f_ASAP7_75t_R register___U14453 ( .A(register__net110028), .Y(register__net90545) );
  BUFx4f_ASAP7_75t_R register___U14454 ( .A(register__net105738), .Y(register__net90541) );
  BUFx4f_ASAP7_75t_R register___U14455 ( .A(register__net103556), .Y(register__net90533) );
  BUFx4f_ASAP7_75t_R register___U14456 ( .A(register__net114109), .Y(register__net90525) );
  BUFx4f_ASAP7_75t_R register___U14457 ( .A(register__net115992), .Y(register__net90521) );
  BUFx4f_ASAP7_75t_R register___U14458 ( .A(register__n9048), .Y(register__n9781) );
  BUFx6f_ASAP7_75t_R register___U14459 ( .A(register__n9783), .Y(register__n9782) );
  BUFx4f_ASAP7_75t_R register___U14460 ( .A(register__n7511), .Y(register__n9783) );
  BUFx6f_ASAP7_75t_R register___U14461 ( .A(register__n9785), .Y(register__n9784) );
  BUFx4f_ASAP7_75t_R register___U14462 ( .A(register__n7798), .Y(register__n9785) );
  BUFx4f_ASAP7_75t_R register___U14463 ( .A(register__n8478), .Y(register__n9787) );
  BUFx6f_ASAP7_75t_R register___U14464 ( .A(register__n9789), .Y(register__n9788) );
  BUFx4f_ASAP7_75t_R register___U14465 ( .A(register__n7196), .Y(register__n9789) );
  BUFx6f_ASAP7_75t_R register___U14466 ( .A(register__n9791), .Y(register__n9790) );
  BUFx4f_ASAP7_75t_R register___U14467 ( .A(register__n7806), .Y(register__n9791) );
  BUFx6f_ASAP7_75t_R register___U14468 ( .A(register__n9793), .Y(register__n9792) );
  BUFx4f_ASAP7_75t_R register___U14469 ( .A(register__n6380), .Y(register__n9793) );
  BUFx6f_ASAP7_75t_R register___U14470 ( .A(register__n9795), .Y(register__n9794) );
  BUFx4f_ASAP7_75t_R register___U14471 ( .A(register__n5885), .Y(register__n9795) );
  BUFx6f_ASAP7_75t_R register___U14472 ( .A(register__n9797), .Y(register__n9796) );
  BUFx4f_ASAP7_75t_R register___U14473 ( .A(register__n8141), .Y(register__n9797) );
  BUFx6f_ASAP7_75t_R register___U14474 ( .A(register__n9799), .Y(register__n9798) );
  BUFx4f_ASAP7_75t_R register___U14475 ( .A(register__n8143), .Y(register__n9799) );
  BUFx6f_ASAP7_75t_R register___U14476 ( .A(register__n9801), .Y(register__n9800) );
  BUFx4f_ASAP7_75t_R register___U14477 ( .A(register__n9051), .Y(register__n9801) );
  BUFx4f_ASAP7_75t_R register___U14478 ( .A(register__n9056), .Y(register__n9803) );
  BUFx6f_ASAP7_75t_R register___U14479 ( .A(register__n9807), .Y(register__n9806) );
  BUFx4f_ASAP7_75t_R register___U14480 ( .A(register__n5209), .Y(register__n9807) );
  BUFx4f_ASAP7_75t_R register___U14481 ( .A(register__net117707), .Y(register__net90453) );
  BUFx6f_ASAP7_75t_R register___U14482 ( .A(register__n9809), .Y(register__n9808) );
  BUFx4f_ASAP7_75t_R register___U14483 ( .A(register__n7518), .Y(register__n9809) );
  BUFx6f_ASAP7_75t_R register___U14484 ( .A(register__n9813), .Y(register__n9812) );
  BUFx4f_ASAP7_75t_R register___U14485 ( .A(register__n7200), .Y(register__n9813) );
  BUFx6f_ASAP7_75t_R register___U14486 ( .A(register__n9815), .Y(register__n9814) );
  BUFx4f_ASAP7_75t_R register___U14487 ( .A(register__n7525), .Y(register__n9815) );
  BUFx6f_ASAP7_75t_R register___U14488 ( .A(register__n9817), .Y(register__n9816) );
  BUFx4f_ASAP7_75t_R register___U14489 ( .A(register__n6937), .Y(register__n9817) );
  BUFx6f_ASAP7_75t_R register___U14490 ( .A(register__n9819), .Y(register__n9818) );
  BUFx4f_ASAP7_75t_R register___U14491 ( .A(register__n7819), .Y(register__n9819) );
  BUFx6f_ASAP7_75t_R register___U14492 ( .A(register__n9821), .Y(register__n9820) );
  BUFx4f_ASAP7_75t_R register___U14493 ( .A(register__n5889), .Y(register__n9821) );
  BUFx6f_ASAP7_75t_R register___U14494 ( .A(register__n9823), .Y(register__n9822) );
  BUFx4f_ASAP7_75t_R register___U14495 ( .A(register__n8158), .Y(register__n9823) );
  BUFx6f_ASAP7_75t_R register___U14496 ( .A(register__n9827), .Y(register__n9826) );
  BUFx4f_ASAP7_75t_R register___U14497 ( .A(register__n6941), .Y(register__n9827) );
  BUFx6f_ASAP7_75t_R register___U14498 ( .A(register__n9829), .Y(register__n9828) );
  BUFx4f_ASAP7_75t_R register___U14499 ( .A(register__n4273), .Y(register__n9829) );
  BUFx4f_ASAP7_75t_R register___U14500 ( .A(register__net103463), .Y(register__net90405) );
  BUFx4f_ASAP7_75t_R register___U14501 ( .A(register__net105686), .Y(register__net90401) );
  BUFx4f_ASAP7_75t_R register___U14502 ( .A(register__net101000), .Y(register__net90397) );
  BUFx4f_ASAP7_75t_R register___U14503 ( .A(register__net105682), .Y(register__net90393) );
  BUFx4f_ASAP7_75t_R register___U14504 ( .A(register__n9077), .Y(register__n9833) );
  BUFx6f_ASAP7_75t_R register___U14505 ( .A(register__n9835), .Y(register__n9834) );
  BUFx4f_ASAP7_75t_R register___U14506 ( .A(register__n7211), .Y(register__n9835) );
  BUFx6f_ASAP7_75t_R register___U14507 ( .A(register__n9839), .Y(register__n9838) );
  BUFx4f_ASAP7_75t_R register___U14508 ( .A(register__n7536), .Y(register__n9839) );
  BUFx4f_ASAP7_75t_R register___U14509 ( .A(register__n9083), .Y(register__n9841) );
  BUFx6f_ASAP7_75t_R register___U14510 ( .A(register__n9844), .Y(register__n9843) );
  BUFx4f_ASAP7_75t_R register___U14511 ( .A(register__n7831), .Y(register__n9844) );
  BUFx6f_ASAP7_75t_R register___U14512 ( .A(register__n9846), .Y(register__n9845) );
  BUFx4f_ASAP7_75t_R register___U14513 ( .A(register__n6122), .Y(register__n9846) );
  BUFx6f_ASAP7_75t_R register___U14514 ( .A(register__n9848), .Y(register__n9847) );
  BUFx4f_ASAP7_75t_R register___U14515 ( .A(register__n3695), .Y(register__n9848) );
  BUFx6f_ASAP7_75t_R register___U14516 ( .A(register__n9850), .Y(register__n9849) );
  BUFx4f_ASAP7_75t_R register___U14517 ( .A(register__n8174), .Y(register__n9850) );
  BUFx6f_ASAP7_75t_R register___U14518 ( .A(register__n9852), .Y(register__n9851) );
  BUFx4f_ASAP7_75t_R register___U14519 ( .A(register__n9092), .Y(register__n9852) );
  BUFx6f_ASAP7_75t_R register___U14520 ( .A(register__n9860), .Y(register__n9859) );
  BUFx4f_ASAP7_75t_R register___U14521 ( .A(register__n7547), .Y(register__n9860) );
  BUFx6f_ASAP7_75t_R register___U14522 ( .A(register__n9864), .Y(register__n9863) );
  BUFx4f_ASAP7_75t_R register___U14523 ( .A(register__n6664), .Y(register__n9864) );
  BUFx6f_ASAP7_75t_R register___U14524 ( .A(register__n9866), .Y(register__n9865) );
  BUFx4f_ASAP7_75t_R register___U14525 ( .A(register__n7552), .Y(register__n9866) );
  BUFx4f_ASAP7_75t_R register___U14526 ( .A(register__n9105), .Y(register__n9868) );
  BUFx6f_ASAP7_75t_R register___U14527 ( .A(register__n9870), .Y(register__n9869) );
  BUFx4f_ASAP7_75t_R register___U14528 ( .A(register__n9108), .Y(register__n9870) );
  BUFx6f_ASAP7_75t_R register___U14529 ( .A(register__n9872), .Y(register__n9871) );
  BUFx4f_ASAP7_75t_R register___U14530 ( .A(register__n4971), .Y(register__n9872) );
  BUFx6f_ASAP7_75t_R register___U14531 ( .A(register__n9874), .Y(register__n9873) );
  BUFx4f_ASAP7_75t_R register___U14532 ( .A(register__n7232), .Y(register__n9874) );
  BUFx6f_ASAP7_75t_R register___U14533 ( .A(register__n9876), .Y(register__n9875) );
  BUFx4f_ASAP7_75t_R register___U14534 ( .A(register__n8191), .Y(register__n9876) );
  BUFx6f_ASAP7_75t_R register___U14535 ( .A(register__n9878), .Y(register__n9877) );
  BUFx4f_ASAP7_75t_R register___U14536 ( .A(register__n8525), .Y(register__n9878) );
  BUFx4f_ASAP7_75t_R register___U14537 ( .A(register__n8530), .Y(register__n9880) );
  BUFx6f_ASAP7_75t_R register___U14538 ( .A(register__n9882), .Y(register__n9881) );
  BUFx4f_ASAP7_75t_R register___U14539 ( .A(register__n5893), .Y(register__n9882) );
  BUFx4f_ASAP7_75t_R register___U14540 ( .A(register__n9122), .Y(register__n9884) );
  BUFx6f_ASAP7_75t_R register___U14541 ( .A(register__n9886), .Y(register__n9885) );
  BUFx4f_ASAP7_75t_R register___U14542 ( .A(register__n8536), .Y(register__n9886) );
  BUFx4f_ASAP7_75t_R register___U14543 ( .A(register__n8195), .Y(register__n9888) );
  BUFx4f_ASAP7_75t_R register___U14544 ( .A(register__n8541), .Y(register__n9890) );
  BUFx4f_ASAP7_75t_R register___U14545 ( .A(register__net109924), .Y(register__net90265) );
  BUFx4f_ASAP7_75t_R register___U14546 ( .A(register__net103364), .Y(register__net90261) );
  BUFx4f_ASAP7_75t_R register___U14547 ( .A(register__net94862), .Y(register__net90258) );
  BUFx4f_ASAP7_75t_R register___U14548 ( .A(register__net107874), .Y(register__net90253) );
  BUFx6f_ASAP7_75t_R register___U14549 ( .A(register__n9892), .Y(register__n9891) );
  BUFx4f_ASAP7_75t_R register___U14550 ( .A(register__n6392), .Y(register__n9892) );
  BUFx6f_ASAP7_75t_R register___U14551 ( .A(register__n9894), .Y(register__n9893) );
  BUFx4f_ASAP7_75t_R register___U14552 ( .A(register__n7571), .Y(register__n9894) );
  BUFx4f_ASAP7_75t_R register___U14553 ( .A(register__net109906), .Y(register__net90237) );
  BUFx4f_ASAP7_75t_R register___U14554 ( .A(register__net105582), .Y(register__net90229) );
  BUFx4f_ASAP7_75t_R register___U14555 ( .A(register__net98210), .Y(register__net90225) );
  BUFx4f_ASAP7_75t_R register___U14556 ( .A(register__net94799), .Y(register__net90221) );
  BUFx4f_ASAP7_75t_R register___U14557 ( .A(register__net98206), .Y(register__net90217) );
  BUFx4f_ASAP7_75t_R register___U14558 ( .A(register__net98201), .Y(register__net90213) );
  BUFx6f_ASAP7_75t_R register___U14559 ( .A(register__n9896), .Y(register__n9895) );
  BUFx4f_ASAP7_75t_R register___U14560 ( .A(register__n7238), .Y(register__n9896) );
  BUFx4f_ASAP7_75t_R register___U14561 ( .A(register__n9141), .Y(register__n9898) );
  BUFx6f_ASAP7_75t_R register___U14562 ( .A(register__n9900), .Y(register__n9899) );
  BUFx4f_ASAP7_75t_R register___U14563 ( .A(register__n8203), .Y(register__n9900) );
  BUFx6f_ASAP7_75t_R register___U14564 ( .A(register__n9904), .Y(register__n9903) );
  BUFx4f_ASAP7_75t_R register___U14565 ( .A(register__n7861), .Y(register__n9904) );
  BUFx6f_ASAP7_75t_R register___U14566 ( .A(register__n9906), .Y(register__n9905) );
  BUFx4f_ASAP7_75t_R register___U14567 ( .A(register__n6677), .Y(register__n9906) );
  BUFx4f_ASAP7_75t_R register___U14568 ( .A(register__n7863), .Y(register__n9908) );
  BUFx4f_ASAP7_75t_R register___U14569 ( .A(register__n9145), .Y(register__n9910) );
  BUFx6f_ASAP7_75t_R register___U14570 ( .A(register__n9912), .Y(register__n9911) );
  BUFx4f_ASAP7_75t_R register___U14571 ( .A(register__n8553), .Y(register__n9912) );
  BUFx6f_ASAP7_75t_R register___U14572 ( .A(register__n9914), .Y(register__n9913) );
  BUFx4f_ASAP7_75t_R register___U14573 ( .A(register__n7240), .Y(register__n9914) );
  BUFx4f_ASAP7_75t_R register___U14574 ( .A(register__net108103), .Y(register__net90169) );
  BUFx6f_ASAP7_75t_R register___U14575 ( .A(register__n9916), .Y(register__n9915) );
  BUFx4f_ASAP7_75t_R register___U14576 ( .A(register__n6080), .Y(register__n9916) );
  BUFx6f_ASAP7_75t_R register___U14577 ( .A(register__n9918), .Y(register__n9917) );
  BUFx4f_ASAP7_75t_R register___U14578 ( .A(register__n5200), .Y(register__n9918) );
  BUFx6f_ASAP7_75t_R register___U14579 ( .A(register__n9920), .Y(register__n9919) );
  BUFx4f_ASAP7_75t_R register___U14580 ( .A(register__n7410), .Y(register__n9920) );
  BUFx6f_ASAP7_75t_R register___U14581 ( .A(register__n9922), .Y(register__n9921) );
  BUFx4f_ASAP7_75t_R register___U14582 ( .A(register__n7412), .Y(register__n9922) );
  BUFx4f_ASAP7_75t_R register___U14583 ( .A(register__net114290), .Y(register__net90149) );
  BUFx4f_ASAP7_75t_R register___U14584 ( .A(register__net108099), .Y(register__net90145) );
  BUFx6f_ASAP7_75t_R register___U14585 ( .A(register__n9924), .Y(register__n9923) );
  BUFx4f_ASAP7_75t_R register___U14586 ( .A(register__n6851), .Y(register__n9924) );
  BUFx6f_ASAP7_75t_R register___U14587 ( .A(register__n9926), .Y(register__n9925) );
  BUFx4f_ASAP7_75t_R register___U14588 ( .A(register__n5861), .Y(register__n9926) );
  BUFx6f_ASAP7_75t_R register___U14589 ( .A(register__n9928), .Y(register__n9927) );
  BUFx4f_ASAP7_75t_R register___U14590 ( .A(register__n7153), .Y(register__n9928) );
  BUFx6f_ASAP7_75t_R register___U14591 ( .A(register__n9930), .Y(register__n9929) );
  BUFx4f_ASAP7_75t_R register___U14592 ( .A(register__n6554), .Y(register__n9930) );
  BUFx6f_ASAP7_75t_R register___U14593 ( .A(register__n9932), .Y(register__n9931) );
  BUFx4f_ASAP7_75t_R register___U14594 ( .A(register__n6317), .Y(register__n9932) );
  BUFx6f_ASAP7_75t_R register___U14595 ( .A(register__n9934), .Y(register__n9933) );
  BUFx4f_ASAP7_75t_R register___U14596 ( .A(register__n7155), .Y(register__n9934) );
  BUFx6f_ASAP7_75t_R register___U14597 ( .A(register__n9936), .Y(register__n9935) );
  BUFx4f_ASAP7_75t_R register___U14598 ( .A(register__n5863), .Y(register__n9936) );
  BUFx4f_ASAP7_75t_R register___U14599 ( .A(register__net101353), .Y(register__net90113) );
  BUFx4f_ASAP7_75t_R register___U14600 ( .A(register__net95646), .Y(register__net90109) );
  BUFx6f_ASAP7_75t_R register___U14601 ( .A(register__n9938), .Y(register__n9937) );
  BUFx4f_ASAP7_75t_R register___U14602 ( .A(register__n7159), .Y(register__n9938) );
  BUFx6f_ASAP7_75t_R register___U14603 ( .A(register__n9940), .Y(register__n9939) );
  BUFx4f_ASAP7_75t_R register___U14604 ( .A(register__n8038), .Y(register__n9940) );
  BUFx6f_ASAP7_75t_R register___U14605 ( .A(register__n9942), .Y(register__n9941) );
  BUFx4f_ASAP7_75t_R register___U14606 ( .A(register__n6556), .Y(register__n9942) );
  BUFx4f_ASAP7_75t_R register___U14607 ( .A(register__net114274), .Y(register__net90093) );
  BUFx6f_ASAP7_75t_R register___U14608 ( .A(register__n9944), .Y(register__n9943) );
  BUFx4f_ASAP7_75t_R register___U14609 ( .A(register__n6558), .Y(register__n9944) );
  BUFx6f_ASAP7_75t_R register___U14610 ( .A(register__n9946), .Y(register__n9945) );
  BUFx4f_ASAP7_75t_R register___U14611 ( .A(register__n3637), .Y(register__n9946) );
  BUFx4f_ASAP7_75t_R register___U14612 ( .A(register__net112503), .Y(register__net90081) );
  BUFx4f_ASAP7_75t_R register___U14613 ( .A(register__net112499), .Y(register__net90077) );
  BUFx6f_ASAP7_75t_R register___U14614 ( .A(register__n9948), .Y(register__n9947) );
  BUFx4f_ASAP7_75t_R register___U14615 ( .A(register__n5526), .Y(register__n9948) );
  BUFx6f_ASAP7_75t_R register___U14616 ( .A(register__n9950), .Y(register__n9949) );
  BUFx4f_ASAP7_75t_R register___U14617 ( .A(register__n8400), .Y(register__n9950) );
  BUFx4f_ASAP7_75t_R register___U14618 ( .A(register__n6853), .Y(register__n9952) );
  BUFx4f_ASAP7_75t_R register___U14619 ( .A(register__net105991), .Y(register__net90061) );
  BUFx6f_ASAP7_75t_R register___U14620 ( .A(register__n9954), .Y(register__n9953) );
  BUFx4f_ASAP7_75t_R register___U14621 ( .A(register__n7414), .Y(register__n9954) );
  BUFx6f_ASAP7_75t_R register___U14622 ( .A(register__n9956), .Y(register__n9955) );
  BUFx4f_ASAP7_75t_R register___U14623 ( .A(register__n7416), .Y(register__n9956) );
  BUFx6f_ASAP7_75t_R register___U14624 ( .A(register__n9958), .Y(register__n9957) );
  BUFx4f_ASAP7_75t_R register___U14625 ( .A(register__n8040), .Y(register__n9958) );
  BUFx6f_ASAP7_75t_R register___U14626 ( .A(register__n9960), .Y(register__n9959) );
  BUFx4f_ASAP7_75t_R register___U14627 ( .A(register__n8042), .Y(register__n9960) );
  BUFx4f_ASAP7_75t_R register___U14628 ( .A(register__net112495), .Y(register__net90041) );
  BUFx4f_ASAP7_75t_R register___U14629 ( .A(register__net110205), .Y(register__net90037) );
  BUFx6f_ASAP7_75t_R register___U14630 ( .A(register__n9964), .Y(register__n9963) );
  BUFx4f_ASAP7_75t_R register___U14631 ( .A(register__n6567), .Y(register__n9964) );
  BUFx6f_ASAP7_75t_R register___U14632 ( .A(register__n9966), .Y(register__n9965) );
  BUFx4f_ASAP7_75t_R register___U14633 ( .A(register__n6324), .Y(register__n9966) );
  BUFx6f_ASAP7_75t_R register___U14634 ( .A(register__n9968), .Y(register__n9967) );
  BUFx4f_ASAP7_75t_R register___U14635 ( .A(register__n6856), .Y(register__n9968) );
  BUFx4f_ASAP7_75t_R register___U14636 ( .A(register__net139226), .Y(register__net90017) );
  BUFx6f_ASAP7_75t_R register___U14637 ( .A(register__n9970), .Y(register__n9969) );
  BUFx4f_ASAP7_75t_R register___U14638 ( .A(register__n7420), .Y(register__n9970) );
  BUFx6f_ASAP7_75t_R register___U14639 ( .A(register__n9972), .Y(register__n9971) );
  BUFx4f_ASAP7_75t_R register___U14640 ( .A(register__n3796), .Y(register__n9972) );
  BUFx6f_ASAP7_75t_R register___U14641 ( .A(register__n9974), .Y(register__n9973) );
  BUFx4f_ASAP7_75t_R register___U14642 ( .A(register__n3798), .Y(register__n9974) );
  BUFx6f_ASAP7_75t_R register___U14643 ( .A(register__n9976), .Y(register__n9975) );
  BUFx4f_ASAP7_75t_R register___U14644 ( .A(register__n7422), .Y(register__n9976) );
  BUFx4f_ASAP7_75t_R register___U14645 ( .A(register__net139206), .Y(register__net89997) );
  BUFx4f_ASAP7_75t_R register___U14646 ( .A(register__net139202), .Y(register__net89993) );
  BUFx6f_ASAP7_75t_R register___U14647 ( .A(register__n9978), .Y(register__n9977) );
  BUFx4f_ASAP7_75t_R register___U14648 ( .A(register__n7424), .Y(register__n9978) );
  BUFx6f_ASAP7_75t_R register___U14649 ( .A(register__n9980), .Y(register__n9979) );
  BUFx4f_ASAP7_75t_R register___U14650 ( .A(register__n7426), .Y(register__n9980) );
  BUFx6f_ASAP7_75t_R register___U14651 ( .A(register__n9982), .Y(register__n9981) );
  BUFx4f_ASAP7_75t_R register___U14652 ( .A(register__n3802), .Y(register__n9982) );
  BUFx6f_ASAP7_75t_R register___U14653 ( .A(register__n9984), .Y(register__n9983) );
  BUFx4f_ASAP7_75t_R register___U14654 ( .A(register__n7428), .Y(register__n9984) );
  BUFx6f_ASAP7_75t_R register___U14655 ( .A(register__n9986), .Y(register__n9985) );
  BUFx4f_ASAP7_75t_R register___U14656 ( .A(register__n3804), .Y(register__n9986) );
  BUFx4f_ASAP7_75t_R register___U14657 ( .A(register__net110197), .Y(register__net89969) );
  BUFx6f_ASAP7_75t_R register___U14658 ( .A(register__n9988), .Y(register__n9987) );
  BUFx4f_ASAP7_75t_R register___U14659 ( .A(register__n6086), .Y(register__n9988) );
  BUFx6f_ASAP7_75t_R register___U14660 ( .A(register__n9990), .Y(register__n9989) );
  BUFx4f_ASAP7_75t_R register___U14661 ( .A(register__n5867), .Y(register__n9990) );
  BUFx6f_ASAP7_75t_R register___U14662 ( .A(register__n9992), .Y(register__n9991) );
  BUFx4f_ASAP7_75t_R register___U14663 ( .A(register__n5869), .Y(register__n9992) );
  BUFx4f_ASAP7_75t_R register___U14664 ( .A(register__net114248), .Y(register__net89953) );
  BUFx6f_ASAP7_75t_R register___U14665 ( .A(register__n9994), .Y(register__n9993) );
  BUFx4f_ASAP7_75t_R register___U14666 ( .A(register__n6330), .Y(register__n9994) );
  BUFx6f_ASAP7_75t_R register___U14667 ( .A(register__n9996), .Y(register__n9995) );
  BUFx4f_ASAP7_75t_R register___U14668 ( .A(register__n5671), .Y(register__n9996) );
  BUFx6f_ASAP7_75t_R register___U14669 ( .A(register__n9998), .Y(register__n9997) );
  BUFx4f_ASAP7_75t_R register___U14670 ( .A(register__n7430), .Y(register__n9998) );
  BUFx6f_ASAP7_75t_R register___U14671 ( .A(register__n10000), .Y(register__n9999) );
  BUFx4f_ASAP7_75t_R register___U14672 ( .A(register__n7447), .Y(register__n10000) );
  BUFx6f_ASAP7_75t_R register___U14673 ( .A(register__n10002), .Y(register__n10001) );
  BUFx4f_ASAP7_75t_R register___U14674 ( .A(register__n8062), .Y(register__n10002) );
  BUFx6f_ASAP7_75t_R register___U14675 ( .A(register__n10005), .Y(register__n10004) );
  BUFx4f_ASAP7_75t_R register___U14676 ( .A(register__n5204), .Y(register__n10005) );
  BUFx6f_ASAP7_75t_R register___U14677 ( .A(register__n10007), .Y(register__n10006) );
  BUFx4f_ASAP7_75t_R register___U14678 ( .A(register__n6868), .Y(register__n10007) );
  BUFx4f_ASAP7_75t_R register___U14679 ( .A(register__n8414), .Y(register__n10009) );
  BUFx4f_ASAP7_75t_R register___U14680 ( .A(register__net98598), .Y(register__net89913) );
  BUFx4f_ASAP7_75t_R register___U14681 ( .A(register__net105913), .Y(register__net89909) );
  BUFx6f_ASAP7_75t_R register___U14682 ( .A(register__n10011), .Y(register__n10010) );
  BUFx4f_ASAP7_75t_R register___U14683 ( .A(register__n8064), .Y(register__n10011) );
  BUFx6f_ASAP7_75t_R register___U14684 ( .A(register__n10015), .Y(register__n10014) );
  BUFx4f_ASAP7_75t_R register___U14685 ( .A(register__n7765), .Y(register__n10015) );
  BUFx6f_ASAP7_75t_R register___U14686 ( .A(register__n10017), .Y(register__n10016) );
  BUFx4f_ASAP7_75t_R register___U14687 ( .A(register__n6579), .Y(register__n10017) );
  BUFx4f_ASAP7_75t_R register___U14688 ( .A(register__net135778), .Y(register__net89889) );
  BUFx6f_ASAP7_75t_R register___U14689 ( .A(register__n10019), .Y(register__n10018) );
  BUFx4f_ASAP7_75t_R register___U14690 ( .A(register__n6581), .Y(register__n10019) );
  BUFx6f_ASAP7_75t_R register___U14691 ( .A(register__n10021), .Y(register__n10020) );
  BUFx4f_ASAP7_75t_R register___U14692 ( .A(register__n6583), .Y(register__n10021) );
  BUFx6f_ASAP7_75t_R register___U14693 ( .A(register__net89878), .Y(register__net89877) );
  BUFx4f_ASAP7_75t_R register___U14694 ( .A(register__net112455), .Y(register__net89878) );
  BUFx6f_ASAP7_75t_R register___U14695 ( .A(register__n10023), .Y(register__n10022) );
  BUFx4f_ASAP7_75t_R register___U14696 ( .A(register__n6585), .Y(register__n10023) );
  BUFx6f_ASAP7_75t_R register___U14697 ( .A(register__n10025), .Y(register__n10024) );
  BUFx4f_ASAP7_75t_R register___U14698 ( .A(register__n6587), .Y(register__n10025) );
  BUFx4f_ASAP7_75t_R register___U14699 ( .A(register__net101273), .Y(register__net89865) );
  BUFx4f_ASAP7_75t_R register___U14700 ( .A(register__net135774), .Y(register__net89861) );
  BUFx6f_ASAP7_75t_R register___U14701 ( .A(register__n10027), .Y(register__n10026) );
  BUFx4f_ASAP7_75t_R register___U14702 ( .A(register__n4039), .Y(register__n10027) );
  BUFx6f_ASAP7_75t_R register___U14703 ( .A(register__n10029), .Y(register__n10028) );
  BUFx4f_ASAP7_75t_R register___U14704 ( .A(register__n4041), .Y(register__n10029) );
  BUFx6f_ASAP7_75t_R register___U14705 ( .A(register__n10031), .Y(register__n10030) );
  BUFx4f_ASAP7_75t_R register___U14706 ( .A(register__n6591), .Y(register__n10031) );
  BUFx4f_ASAP7_75t_R register___U14707 ( .A(register__net95571), .Y(register__net89846) );
  BUFx4f_ASAP7_75t_R register___U14708 ( .A(register__n8889), .Y(register__n10035) );
  BUFx3_ASAP7_75t_R register___U14709 ( .A(register__n8838), .Y(register__n10037) );
  BUFx6f_ASAP7_75t_R register___U14710 ( .A(register__n10043), .Y(register__n10042) );
  BUFx4f_ASAP7_75t_R register___U14711 ( .A(register__n8070), .Y(register__n10043) );
  BUFx4f_ASAP7_75t_R register___U14712 ( .A(register__net95557), .Y(register__net89814) );
  BUFx4f_ASAP7_75t_R register___U14713 ( .A(register__n8892), .Y(register__n10045) );
  BUFx4f_ASAP7_75t_R register___U14714 ( .A(register__n8899), .Y(register__n10051) );
  BUFx4f_ASAP7_75t_R register___U14715 ( .A(register__net98553), .Y(register__net89794) );
  BUFx6f_ASAP7_75t_R register___U14716 ( .A(register__n10053), .Y(register__n10052) );
  BUFx4f_ASAP7_75t_R register___U14717 ( .A(register__n7453), .Y(register__n10053) );
  BUFx6f_ASAP7_75t_R register___U14718 ( .A(register__n10055), .Y(register__n10054) );
  BUFx4f_ASAP7_75t_R register___U14719 ( .A(register__n7455), .Y(register__n10055) );
  BUFx6f_ASAP7_75t_R register___U14720 ( .A(register__n10057), .Y(register__n10056) );
  BUFx4f_ASAP7_75t_R register___U14721 ( .A(register__n5673), .Y(register__n10057) );
  BUFx4f_ASAP7_75t_R register___U14722 ( .A(register__net105883), .Y(register__net89777) );
  BUFx4f_ASAP7_75t_R register___U14723 ( .A(register__net105879), .Y(register__net89773) );
  BUFx6f_ASAP7_75t_R register___U14724 ( .A(register__n10059), .Y(register__n10058) );
  BUFx4f_ASAP7_75t_R register___U14725 ( .A(register__n7460), .Y(register__n10059) );
  BUFx6f_ASAP7_75t_R register___U14726 ( .A(register__n10061), .Y(register__n10060) );
  BUFx4f_ASAP7_75t_R register___U14727 ( .A(register__n7462), .Y(register__n10061) );
  BUFx6f_ASAP7_75t_R register___U14728 ( .A(register__n10063), .Y(register__n10062) );
  BUFx4f_ASAP7_75t_R register___U14729 ( .A(register__n8076), .Y(register__n10063) );
  BUFx6f_ASAP7_75t_R register___U14730 ( .A(register__n10065), .Y(register__n10064) );
  BUFx4f_ASAP7_75t_R register___U14731 ( .A(register__n8943), .Y(register__n10065) );
  BUFx6f_ASAP7_75t_R register___U14732 ( .A(register__n10067), .Y(register__n10066) );
  BUFx4f_ASAP7_75t_R register___U14733 ( .A(register__n8078), .Y(register__n10067) );
  BUFx6f_ASAP7_75t_R register___U14734 ( .A(register__n10069), .Y(register__n10068) );
  BUFx4f_ASAP7_75t_R register___U14735 ( .A(register__n8948), .Y(register__n10069) );
  BUFx6f_ASAP7_75t_R register___U14736 ( .A(register__n10071), .Y(register__n10070) );
  BUFx4f_ASAP7_75t_R register___U14737 ( .A(register__n7475), .Y(register__n10071) );
  BUFx4f_ASAP7_75t_R register___U14738 ( .A(register__net98542), .Y(register__net89742) );
  BUFx4f_ASAP7_75t_R register___U14739 ( .A(register__n8950), .Y(register__n10073) );
  BUFx6f_ASAP7_75t_R register___U14740 ( .A(register__n10077), .Y(register__n10076) );
  BUFx4f_ASAP7_75t_R register___U14741 ( .A(register__n7769), .Y(register__n10077) );
  BUFx4f_ASAP7_75t_R register___U14742 ( .A(register__n8956), .Y(register__n10079) );
  BUFx4f_ASAP7_75t_R register___U14743 ( .A(register__n8959), .Y(register__n10081) );
  BUFx4f_ASAP7_75t_R register___U14744 ( .A(register__net103641), .Y(register__net89717) );
  BUFx4f_ASAP7_75t_R register___U14745 ( .A(register__net95372), .Y(register__net89714) );
  BUFx6f_ASAP7_75t_R register___U14746 ( .A(register__n10083), .Y(register__n10082) );
  BUFx4f_ASAP7_75t_R register___U14747 ( .A(register__n8080), .Y(register__n10083) );
  BUFx6f_ASAP7_75t_R register___U14748 ( .A(register__n10085), .Y(register__n10084) );
  BUFx4f_ASAP7_75t_R register___U14749 ( .A(register__n7482), .Y(register__n10085) );
  BUFx6f_ASAP7_75t_R register___U14750 ( .A(register__n10087), .Y(register__n10086) );
  BUFx4f_ASAP7_75t_R register___U14751 ( .A(register__n7484), .Y(register__n10087) );
  BUFx6f_ASAP7_75t_R register___U14752 ( .A(register__n10089), .Y(register__n10088) );
  BUFx4f_ASAP7_75t_R register___U14753 ( .A(register__n8085), .Y(register__n10089) );
  BUFx4f_ASAP7_75t_R register___U14754 ( .A(register__net103630), .Y(register__net89689) );
  BUFx4f_ASAP7_75t_R register___U14755 ( .A(register__net95365), .Y(register__net89686) );
  BUFx6f_ASAP7_75t_R register___U14756 ( .A(register__n10092), .Y(register__n10091) );
  BUFx4f_ASAP7_75t_R register___U14757 ( .A(register__n7773), .Y(register__n10092) );
  BUFx4f_ASAP7_75t_R register___U14758 ( .A(register__net95321), .Y(register__net89662) );
  BUFx4f_ASAP7_75t_R register___U14759 ( .A(register__net95310), .Y(register__net89658) );
  BUFx6f_ASAP7_75t_R register___U14760 ( .A(register__n10099), .Y(register__n10098) );
  BUFx4f_ASAP7_75t_R register___U14761 ( .A(register__n3806), .Y(register__n10099) );
  BUFx4f_ASAP7_75t_R register___U14762 ( .A(register__net112427), .Y(register__net89649) );
  BUFx4f_ASAP7_75t_R register___U14763 ( .A(register__net114196), .Y(register__net89641) );
  BUFx6f_ASAP7_75t_R register___U14764 ( .A(register__n10103), .Y(register__n10102) );
  BUFx4f_ASAP7_75t_R register___U14765 ( .A(register__n7775), .Y(register__n10103) );
  BUFx6f_ASAP7_75t_R register___U14766 ( .A(register__n10105), .Y(register__n10104) );
  BUFx4f_ASAP7_75t_R register___U14767 ( .A(register__n6346), .Y(register__n10105) );
  BUFx6f_ASAP7_75t_R register___U14768 ( .A(register__n10107), .Y(register__n10106) );
  BUFx4f_ASAP7_75t_R register___U14769 ( .A(register__n6874), .Y(register__n10107) );
  BUFx4f_ASAP7_75t_R register___U14770 ( .A(register__net127331), .Y(register__net89617) );
  BUFx4f_ASAP7_75t_R register___U14771 ( .A(register__net139186), .Y(register__net89613) );
  BUFx6f_ASAP7_75t_R register___U14772 ( .A(register__n10111), .Y(register__n10110) );
  BUFx4f_ASAP7_75t_R register___U14773 ( .A(register__n6601), .Y(register__n10111) );
  BUFx6f_ASAP7_75t_R register___U14774 ( .A(register__n10113), .Y(register__n10112) );
  BUFx4f_ASAP7_75t_R register___U14775 ( .A(register__n6352), .Y(register__n10113) );
  BUFx4f_ASAP7_75t_R register___U14776 ( .A(register__net98508), .Y(register__net89601) );
  BUFx4f_ASAP7_75t_R register___U14777 ( .A(register__net95227), .Y(register__net89598) );
  BUFx4f_ASAP7_75t_R register___U14778 ( .A(register__net108010), .Y(register__net89594) );
  BUFx4f_ASAP7_75t_R register___U14779 ( .A(register__net103611), .Y(register__net89590) );
  BUFx4f_ASAP7_75t_R register___U14780 ( .A(register__net95220), .Y(register__net89582) );
  BUFx6f_ASAP7_75t_R register___U14781 ( .A(register__n10115), .Y(register__n10114) );
  BUFx4f_ASAP7_75t_R register___U14782 ( .A(register__n7183), .Y(register__n10115) );
  BUFx6f_ASAP7_75t_R register___U14783 ( .A(register__n10117), .Y(register__n10116) );
  BUFx4f_ASAP7_75t_R register___U14784 ( .A(register__n6881), .Y(register__n10117) );
  BUFx6f_ASAP7_75t_R register___U14785 ( .A(register__n10119), .Y(register__n10118) );
  BUFx4f_ASAP7_75t_R register___U14786 ( .A(register__n6356), .Y(register__n10119) );
  BUFx4f_ASAP7_75t_R register___U14787 ( .A(register__n6364), .Y(register__n10125) );
  BUFx6f_ASAP7_75t_R register___U14788 ( .A(register__n10127), .Y(register__n10126) );
  BUFx4f_ASAP7_75t_R register___U14789 ( .A(register__n7783), .Y(register__n10127) );
  BUFx6f_ASAP7_75t_R register___U14790 ( .A(register__n10131), .Y(register__n10130) );
  BUFx4f_ASAP7_75t_R register___U14791 ( .A(register__n6607), .Y(register__n10131) );
  BUFx4f_ASAP7_75t_R register___U14792 ( .A(register__n8445), .Y(register__n10133) );
  BUFx6f_ASAP7_75t_R register___U14793 ( .A(register__n10135), .Y(register__n10134) );
  BUFx4f_ASAP7_75t_R register___U14794 ( .A(register__n6109), .Y(register__n10135) );
  BUFx3_ASAP7_75t_R register___U14795 ( .A(register__n8843), .Y(register__n10141) );
  BUFx6f_ASAP7_75t_R register___U14796 ( .A(register__n10143), .Y(register__n10142) );
  BUFx4f_ASAP7_75t_R register___U14797 ( .A(register__n6888), .Y(register__n10143) );
  BUFx6f_ASAP7_75t_R register___U14798 ( .A(register__n10145), .Y(register__n10144) );
  BUFx4f_ASAP7_75t_R register___U14799 ( .A(register__n6367), .Y(register__n10145) );
  BUFx6f_ASAP7_75t_R register___U14800 ( .A(register__n10147), .Y(register__n10146) );
  BUFx4f_ASAP7_75t_R register___U14801 ( .A(register__n8113), .Y(register__n10147) );
  BUFx4f_ASAP7_75t_R register___U14802 ( .A(register__n8118), .Y(register__n10149) );
  BUFx6f_ASAP7_75t_R register___U14803 ( .A(register__n10151), .Y(register__n10150) );
  BUFx4f_ASAP7_75t_R register___U14804 ( .A(register__n8452), .Y(register__n10151) );
  BUFx4f_ASAP7_75t_R register___U14805 ( .A(register__n9019), .Y(register__n10156) );
  BUFx4f_ASAP7_75t_R register___U14806 ( .A(register__n9024), .Y(register__n10161) );
  BUFx6f_ASAP7_75t_R register___U14807 ( .A(register__n10163), .Y(register__n10162) );
  BUFx4f_ASAP7_75t_R register___U14808 ( .A(register__n6114), .Y(register__n10163) );
  BUFx4f_ASAP7_75t_R register___U14809 ( .A(register__net112381), .Y(register__net89461) );
  BUFx6f_ASAP7_75t_R register___U14810 ( .A(register__n10168), .Y(register__n10167) );
  BUFx4f_ASAP7_75t_R register___U14811 ( .A(register__n6917), .Y(register__n10168) );
  BUFx6f_ASAP7_75t_R register___U14812 ( .A(register__n10170), .Y(register__n10169) );
  BUFx4f_ASAP7_75t_R register___U14813 ( .A(register__n6919), .Y(register__n10170) );
  BUFx6f_ASAP7_75t_R register___U14814 ( .A(register__n10172), .Y(register__n10171) );
  BUFx4f_ASAP7_75t_R register___U14815 ( .A(register__n6373), .Y(register__n10172) );
  BUFx6f_ASAP7_75t_R register___U14816 ( .A(register__n10174), .Y(register__n10173) );
  BUFx4f_ASAP7_75t_R register___U14817 ( .A(register__n5875), .Y(register__n10174) );
  BUFx4f_ASAP7_75t_R register___U14818 ( .A(register__n9043), .Y(register__n10176) );
  BUFx4f_ASAP7_75t_R register___U14819 ( .A(register__net112343), .Y(register__net89425) );
  BUFx4f_ASAP7_75t_R register___U14820 ( .A(register__net105734), .Y(register__net89421) );
  BUFx4f_ASAP7_75t_R register___U14821 ( .A(register__net103566), .Y(register__net89417) );
  BUFx4f_ASAP7_75t_R register___U14822 ( .A(register__net112339), .Y(register__net89413) );
  BUFx4f_ASAP7_75t_R register___U14823 ( .A(register__net135762), .Y(register__net89409) );
  BUFx4f_ASAP7_75t_R register___U14824 ( .A(register__net98400), .Y(register__net89406) );
  BUFx4f_ASAP7_75t_R register___U14825 ( .A(register__net119326), .Y(register__net89401) );
  BUFx4f_ASAP7_75t_R register___U14826 ( .A(register__net139178), .Y(register__net89397) );
  BUFx4f_ASAP7_75t_R register___U14827 ( .A(register__net115996), .Y(register__net89393) );
  BUFx4f_ASAP7_75t_R register___U14828 ( .A(register__net95063), .Y(register__net89390) );
  BUFx6f_ASAP7_75t_R register___U14829 ( .A(register__n10178), .Y(register__n10177) );
  BUFx4f_ASAP7_75t_R register___U14830 ( .A(register__n6627), .Y(register__n10178) );
  BUFx6f_ASAP7_75t_R register___U14831 ( .A(register__n10180), .Y(register__n10179) );
  BUFx4f_ASAP7_75t_R register___U14832 ( .A(register__n8130), .Y(register__n10180) );
  BUFx6f_ASAP7_75t_R register___U14833 ( .A(register__n10182), .Y(register__n10181) );
  BUFx4f_ASAP7_75t_R register___U14834 ( .A(register__n8135), .Y(register__n10182) );
  BUFx6f_ASAP7_75t_R register___U14835 ( .A(register__n10184), .Y(register__n10183) );
  BUFx4f_ASAP7_75t_R register___U14836 ( .A(register__n3808), .Y(register__n10184) );
  BUFx6f_ASAP7_75t_R register___U14837 ( .A(register__n10186), .Y(register__n10185) );
  BUFx4f_ASAP7_75t_R register___U14838 ( .A(register__n6632), .Y(register__n10186) );
  BUFx6f_ASAP7_75t_R register___U14839 ( .A(register__n10190), .Y(register__n10189) );
  BUFx4f_ASAP7_75t_R register___U14840 ( .A(register__n5677), .Y(register__n10190) );
  BUFx6f_ASAP7_75t_R register___U14841 ( .A(register__n10192), .Y(register__n10191) );
  BUFx4f_ASAP7_75t_R register___U14842 ( .A(register__n5879), .Y(register__n10192) );
  BUFx6f_ASAP7_75t_R register___U14843 ( .A(register__n10194), .Y(register__n10193) );
  BUFx4f_ASAP7_75t_R register___U14844 ( .A(register__n5881), .Y(register__n10194) );
  BUFx6f_ASAP7_75t_R register___U14845 ( .A(register__n10196), .Y(register__n10195) );
  BUFx4f_ASAP7_75t_R register___U14846 ( .A(register__n5883), .Y(register__n10196) );
  BUFx6f_ASAP7_75t_R register___U14847 ( .A(register__n10198), .Y(register__n10197) );
  BUFx4f_ASAP7_75t_R register___U14848 ( .A(register__n6634), .Y(register__n10198) );
  BUFx6f_ASAP7_75t_R register___U14849 ( .A(register__n10200), .Y(register__n10199) );
  BUFx4f_ASAP7_75t_R register___U14850 ( .A(register__n7516), .Y(register__n10200) );
  BUFx6f_ASAP7_75t_R register___U14851 ( .A(register__n10202), .Y(register__n10201) );
  BUFx4f_ASAP7_75t_R register___U14852 ( .A(register__n4124), .Y(register__n10202) );
  BUFx4f_ASAP7_75t_R register___U14853 ( .A(register__n8486), .Y(register__n10204) );
  BUFx6f_ASAP7_75t_R register___U14854 ( .A(register__n10207), .Y(register__n10206) );
  BUFx4f_ASAP7_75t_R register___U14855 ( .A(register__n6636), .Y(register__n10207) );
  BUFx6f_ASAP7_75t_R register___U14856 ( .A(register__n10209), .Y(register__n10208) );
  BUFx4f_ASAP7_75t_R register___U14857 ( .A(register__n6382), .Y(register__n10209) );
  BUFx6f_ASAP7_75t_R register___U14858 ( .A(register__n10211), .Y(register__n10210) );
  BUFx4f_ASAP7_75t_R register___U14859 ( .A(register__n3810), .Y(register__n10211) );
  BUFx6f_ASAP7_75t_R register___U14860 ( .A(register__n10213), .Y(register__n10212) );
  BUFx4f_ASAP7_75t_R register___U14861 ( .A(register__n6928), .Y(register__n10213) );
  BUFx6f_ASAP7_75t_R register___U14862 ( .A(register__n10215), .Y(register__n10214) );
  BUFx4f_ASAP7_75t_R register___U14863 ( .A(register__n6933), .Y(register__n10215) );
  BUFx6f_ASAP7_75t_R register___U14864 ( .A(register__n10217), .Y(register__n10216) );
  BUFx4f_ASAP7_75t_R register___U14865 ( .A(register__n6638), .Y(register__n10217) );
  BUFx6f_ASAP7_75t_R register___U14866 ( .A(register__n10220), .Y(register__n10219) );
  BUFx4f_ASAP7_75t_R register___U14867 ( .A(register__n9059), .Y(register__n10220) );
  BUFx6f_ASAP7_75t_R register___U14868 ( .A(register__n10222), .Y(register__n10221) );
  BUFx4f_ASAP7_75t_R register___U14869 ( .A(register__n8488), .Y(register__n10222) );
  BUFx4f_ASAP7_75t_R register___U14870 ( .A(register__net101045), .Y(register__net89289) );
  BUFx4f_ASAP7_75t_R register___U14871 ( .A(register__net101038), .Y(register__net89286) );
  BUFx4f_ASAP7_75t_R register___U14872 ( .A(register__net112295), .Y(register__net89281) );
  BUFx4f_ASAP7_75t_R register___U14873 ( .A(register__net107970), .Y(register__net89277) );
  BUFx4f_ASAP7_75t_R register___U14874 ( .A(register__net115974), .Y(register__net89273) );
  BUFx6f_ASAP7_75t_R register___U14875 ( .A(register__n10226), .Y(register__n10225) );
  BUFx4f_ASAP7_75t_R register___U14876 ( .A(register__n8153), .Y(register__n10226) );
  BUFx6f_ASAP7_75t_R register___U14877 ( .A(register__n10228), .Y(register__n10227) );
  BUFx4f_ASAP7_75t_R register___U14878 ( .A(register__n7202), .Y(register__n10228) );
  BUFx6f_ASAP7_75t_R register___U14879 ( .A(register__n10230), .Y(register__n10229) );
  BUFx4f_ASAP7_75t_R register___U14880 ( .A(register__n6939), .Y(register__n10230) );
  BUFx6f_ASAP7_75t_R register___U14881 ( .A(register__n10232), .Y(register__n10231) );
  BUFx4f_ASAP7_75t_R register___U14882 ( .A(register__n7527), .Y(register__n10232) );
  BUFx4f_ASAP7_75t_R register___U14883 ( .A(register__n8499), .Y(register__n10234) );
  BUFx4f_ASAP7_75t_R register___U14884 ( .A(register__n9074), .Y(register__n10236) );
  BUFx6f_ASAP7_75t_R register___U14885 ( .A(register__n10238), .Y(register__n10237) );
  BUFx4f_ASAP7_75t_R register___U14886 ( .A(register__n5682), .Y(register__n10238) );
  BUFx6f_ASAP7_75t_R register___U14887 ( .A(register__n10240), .Y(register__n10239) );
  BUFx4f_ASAP7_75t_R register___U14888 ( .A(register__n7204), .Y(register__n10240) );
  BUFx6f_ASAP7_75t_R register___U14889 ( .A(register__n10242), .Y(register__n10241) );
  BUFx4f_ASAP7_75t_R register___U14890 ( .A(register__n8163), .Y(register__n10242) );
  BUFx6f_ASAP7_75t_R register___U14891 ( .A(register__n10244), .Y(register__n10243) );
  BUFx4f_ASAP7_75t_R register___U14892 ( .A(register__n4479), .Y(register__n10244) );
  BUFx6f_ASAP7_75t_R register___U14893 ( .A(register__n10246), .Y(register__n10245) );
  BUFx4f_ASAP7_75t_R register___U14894 ( .A(register__n7206), .Y(register__n10246) );
  BUFx6f_ASAP7_75t_R register___U14895 ( .A(register__n10248), .Y(register__n10247) );
  BUFx4f_ASAP7_75t_R register___U14896 ( .A(register__n8502), .Y(register__n10248) );
  BUFx6f_ASAP7_75t_R register___U14897 ( .A(register__n10250), .Y(register__n10249) );
  BUFx4f_ASAP7_75t_R register___U14898 ( .A(register__n6946), .Y(register__n10250) );
  BUFx4f_ASAP7_75t_R register___U14899 ( .A(register__net100990), .Y(register__net89213) );
  BUFx4f_ASAP7_75t_R register___U14900 ( .A(register__net94980), .Y(register__net89210) );
  BUFx4f_ASAP7_75t_R register___U14901 ( .A(register__net103453), .Y(register__net89205) );
  BUFx6f_ASAP7_75t_R register___U14902 ( .A(register__n10252), .Y(register__n10251) );
  BUFx4f_ASAP7_75t_R register___U14903 ( .A(register__n6642), .Y(register__n10252) );
  BUFx4f_ASAP7_75t_R register___U14904 ( .A(register__n7826), .Y(register__n10254) );
  BUFx6f_ASAP7_75t_R register___U14905 ( .A(register__n10256), .Y(register__n10255) );
  BUFx4f_ASAP7_75t_R register___U14906 ( .A(register__n7213), .Y(register__n10256) );
  BUFx6f_ASAP7_75t_R register___U14907 ( .A(register__n10258), .Y(register__n10257) );
  BUFx4f_ASAP7_75t_R register___U14908 ( .A(register__n3814), .Y(register__n10258) );
  BUFx6f_ASAP7_75t_R register___U14909 ( .A(register__n10260), .Y(register__n10259) );
  BUFx4f_ASAP7_75t_R register___U14910 ( .A(register__n6647), .Y(register__n10260) );
  BUFx4f_ASAP7_75t_R register___U14911 ( .A(register__n9080), .Y(register__n10262) );
  BUFx6f_ASAP7_75t_R register___U14912 ( .A(register__n10264), .Y(register__n10263) );
  BUFx4f_ASAP7_75t_R register___U14913 ( .A(register__n6120), .Y(register__n10264) );
  BUFx6f_ASAP7_75t_R register___U14914 ( .A(register__n10266), .Y(register__n10265) );
  BUFx4f_ASAP7_75t_R register___U14915 ( .A(register__n8167), .Y(register__n10266) );
  BUFx6f_ASAP7_75t_R register___U14916 ( .A(register__n10270), .Y(register__n10269) );
  BUFx4f_ASAP7_75t_R register___U14917 ( .A(register__n8507), .Y(register__n10270) );
  BUFx4f_ASAP7_75t_R register___U14918 ( .A(register__n9086), .Y(register__n10272) );
  BUFx4f_ASAP7_75t_R register___U14919 ( .A(register__n8176), .Y(register__n10274) );
  BUFx4f_ASAP7_75t_R register___U14920 ( .A(register__n9089), .Y(register__n10276) );
  BUFx6f_ASAP7_75t_R register___U14921 ( .A(register__n10278), .Y(register__n10277) );
  BUFx4f_ASAP7_75t_R register___U14922 ( .A(register__n7227), .Y(register__n10278) );
  BUFx6f_ASAP7_75t_R register___U14923 ( .A(register__n10280), .Y(register__n10279) );
  BUFx4f_ASAP7_75t_R register___U14924 ( .A(register__n6659), .Y(register__n10280) );
  BUFx4f_ASAP7_75t_R register___U14925 ( .A(register__n8184), .Y(register__n10282) );
  BUFx6f_ASAP7_75t_R register___U14926 ( .A(register__n10284), .Y(register__n10283) );
  BUFx4f_ASAP7_75t_R register___U14927 ( .A(register__n7545), .Y(register__n10284) );
  BUFx6f_ASAP7_75t_R register___U14928 ( .A(register__n10286), .Y(register__n10285) );
  BUFx4f_ASAP7_75t_R register___U14929 ( .A(register__n3816), .Y(register__n10286) );
  BUFx6f_ASAP7_75t_R register___U14930 ( .A(register__n10288), .Y(register__n10287) );
  BUFx4f_ASAP7_75t_R register___U14931 ( .A(register__n7837), .Y(register__n10288) );
  BUFx4f_ASAP7_75t_R register___U14932 ( .A(register__n9097), .Y(register__n10290) );
  BUFx6f_ASAP7_75t_R register___U14933 ( .A(register__n10294), .Y(register__n10293) );
  BUFx4f_ASAP7_75t_R register___U14934 ( .A(register__n7839), .Y(register__n10294) );
  BUFx4f_ASAP7_75t_R register___U14935 ( .A(register__n8517), .Y(register__n10296) );
  BUFx6f_ASAP7_75t_R register___U14936 ( .A(register__n10298), .Y(register__n10297) );
  BUFx4f_ASAP7_75t_R register___U14937 ( .A(register__n5891), .Y(register__n10298) );
  BUFx6f_ASAP7_75t_R register___U14938 ( .A(register__n10300), .Y(register__n10299) );
  BUFx4f_ASAP7_75t_R register___U14939 ( .A(register__n8520), .Y(register__n10300) );
  BUFx4f_ASAP7_75t_R register___U14940 ( .A(register__n9113), .Y(register__n10302) );
  BUFx4f_ASAP7_75t_R register___U14941 ( .A(register__n9116), .Y(register__n10304) );
  BUFx4f_ASAP7_75t_R register___U14942 ( .A(register__n9119), .Y(register__n10306) );
  BUFx6f_ASAP7_75t_R register___U14943 ( .A(register__n10308), .Y(register__n10307) );
  BUFx4f_ASAP7_75t_R register___U14944 ( .A(register__n4043), .Y(register__n10308) );
  BUFx6f_ASAP7_75t_R register___U14945 ( .A(register__n10310), .Y(register__n10309) );
  BUFx4f_ASAP7_75t_R register___U14946 ( .A(register__n7559), .Y(register__n10310) );
  BUFx6f_ASAP7_75t_R register___U14947 ( .A(register__n10312), .Y(register__n10311) );
  BUFx4f_ASAP7_75t_R register___U14948 ( .A(register__n3818), .Y(register__n10312) );
  BUFx6f_ASAP7_75t_R register___U14949 ( .A(register__n10316), .Y(register__n10315) );
  BUFx4f_ASAP7_75t_R register___U14950 ( .A(register__n6388), .Y(register__n10316) );
  BUFx6f_ASAP7_75t_R register___U14951 ( .A(register__n10320), .Y(register__n10319) );
  BUFx4f_ASAP7_75t_R register___U14952 ( .A(register__n7236), .Y(register__n10320) );
  BUFx6f_ASAP7_75t_R register___U14953 ( .A(register__n10322), .Y(register__n10321) );
  BUFx4f_ASAP7_75t_R register___U14954 ( .A(register__n6967), .Y(register__n10322) );
  BUFx4f_ASAP7_75t_R register___U14955 ( .A(register__net100892), .Y(register__net89053) );
  BUFx4f_ASAP7_75t_R register___U14956 ( .A(register__net100885), .Y(register__net89050) );
  BUFx4f_ASAP7_75t_R register___U14957 ( .A(register__net98224), .Y(register__net89046) );
  BUFx4f_ASAP7_75t_R register___U14958 ( .A(register__net107866), .Y(register__net89037) );
  BUFx6f_ASAP7_75t_R register___U14959 ( .A(register__n10324), .Y(register__n10323) );
  BUFx4f_ASAP7_75t_R register___U14960 ( .A(register__n6969), .Y(register__n10324) );
  BUFx6f_ASAP7_75t_R register___U14961 ( .A(register__n10326), .Y(register__n10325) );
  BUFx4f_ASAP7_75t_R register___U14962 ( .A(register__n6673), .Y(register__n10326) );
  BUFx4f_ASAP7_75t_R register___U14963 ( .A(register__n9125), .Y(register__n10328) );
  BUFx6f_ASAP7_75t_R register___U14964 ( .A(register__n10330), .Y(register__n10329) );
  BUFx4f_ASAP7_75t_R register___U14965 ( .A(register__n9128), .Y(register__n10330) );
  BUFx4f_ASAP7_75t_R register___U14966 ( .A(register__net98191), .Y(register__net89017) );
  BUFx4f_ASAP7_75t_R register___U14967 ( .A(register__net94795), .Y(register__net89005) );
  BUFx4f_ASAP7_75t_R register___U14968 ( .A(register__net98184), .Y(register__net89002) );
  BUFx4f_ASAP7_75t_R register___U14969 ( .A(register__net94785), .Y(register__net88997) );
  BUFx6f_ASAP7_75t_R register___U14970 ( .A(register__n10332), .Y(register__n10331) );
  BUFx4f_ASAP7_75t_R register___U14971 ( .A(register__n8546), .Y(register__n10332) );
  BUFx4f_ASAP7_75t_R register___U14972 ( .A(register__n8551), .Y(register__n10334) );
  BUFx4f_ASAP7_75t_R register___U14973 ( .A(register__n9143), .Y(register__n10336) );
  BUFx6f_ASAP7_75t_R register___U14974 ( .A(register__n10338), .Y(register__n10337) );
  BUFx4f_ASAP7_75t_R register___U14975 ( .A(register__n8208), .Y(register__n10338) );
  BUFx6f_ASAP7_75t_R register___U14976 ( .A(register__net88978), .Y(register__net88977) );
  BUFx4f_ASAP7_75t_R register___U14977 ( .A(register__net95678), .Y(register__net88978) );
  BUFx6f_ASAP7_75t_R register___U14978 ( .A(register__n10340), .Y(register__n10339) );
  BUFx4f_ASAP7_75t_R register___U14979 ( .A(register__n8857), .Y(register__n10340) );
  BUFx6f_ASAP7_75t_R register___U14980 ( .A(register__n10342), .Y(register__n10341) );
  BUFx4f_ASAP7_75t_R register___U14981 ( .A(register__n8883), .Y(register__n10342) );
  BUFx6f_ASAP7_75t_R register___U14982 ( .A(register__n10344), .Y(register__n10343) );
  BUFx4f_ASAP7_75t_R register___U14983 ( .A(register__n8885), .Y(register__n10344) );
  BUFx6f_ASAP7_75t_R register___U14984 ( .A(register__n10346), .Y(register__n10345) );
  BUFx4f_ASAP7_75t_R register___U14985 ( .A(register__n8406), .Y(register__n10346) );
  BUFx6f_ASAP7_75t_R register___U14986 ( .A(register__net88958), .Y(register__net88957) );
  BUFx4f_ASAP7_75t_R register___U14987 ( .A(register__net105909), .Y(register__net88958) );
  BUFx6f_ASAP7_75t_R register___U14988 ( .A(register__n10348), .Y(register__n10347) );
  BUFx4f_ASAP7_75t_R register___U14989 ( .A(register__n6870), .Y(register__n10348) );
  BUFx6f_ASAP7_75t_R register___U14990 ( .A(register__net88950), .Y(register__net88949) );
  BUFx4f_ASAP7_75t_R register___U14991 ( .A(register__net98578), .Y(register__net88950) );
  BUFx6f_ASAP7_75t_R register___U14992 ( .A(register__n10350), .Y(register__n10349) );
  BUFx4f_ASAP7_75t_R register___U14993 ( .A(register__n7449), .Y(register__n10350) );
  BUFx6f_ASAP7_75t_R register___U14994 ( .A(register__n10352), .Y(register__n10351) );
  BUFx4f_ASAP7_75t_R register___U14995 ( .A(register__n7767), .Y(register__n10352) );
  BUFx6f_ASAP7_75t_R register___U14996 ( .A(register__n10354), .Y(register__n10353) );
  BUFx4f_ASAP7_75t_R register___U14997 ( .A(register__n8072), .Y(register__n10354) );
  BUFx6f_ASAP7_75t_R register___U14998 ( .A(register__n10358), .Y(register__n10357) );
  BUFx4f_ASAP7_75t_R register___U14999 ( .A(register__n8941), .Y(register__n10358) );
  BUFx6f_ASAP7_75t_R register___U15000 ( .A(register__n10360), .Y(register__n10359) );
  BUFx4f_ASAP7_75t_R register___U15001 ( .A(register__n8429), .Y(register__n10360) );
  BUFx6f_ASAP7_75t_R register___U15002 ( .A(register__n10362), .Y(register__n10361) );
  BUFx4f_ASAP7_75t_R register___U15003 ( .A(register__n8074), .Y(register__n10362) );
  BUFx6f_ASAP7_75t_R register___U15004 ( .A(register__n10364), .Y(register__n10363) );
  BUFx4f_ASAP7_75t_R register___U15005 ( .A(register__n8431), .Y(register__n10364) );
  BUFx4f_ASAP7_75t_R register___U15006 ( .A(register__net108035), .Y(register__net88913) );
  BUFx6f_ASAP7_75t_R register___U15007 ( .A(register__n10366), .Y(register__n10365) );
  BUFx4f_ASAP7_75t_R register___U15008 ( .A(register__n7179), .Y(register__n10366) );
  BUFx6f_ASAP7_75t_R register___U15009 ( .A(register__n10368), .Y(register__n10367) );
  BUFx4f_ASAP7_75t_R register___U15010 ( .A(register__n7469), .Y(register__n10368) );
  BUFx6f_ASAP7_75t_R register___U15011 ( .A(register__n10370), .Y(register__n10369) );
  BUFx4f_ASAP7_75t_R register___U15012 ( .A(register__n7471), .Y(register__n10370) );
  BUFx6f_ASAP7_75t_R register___U15013 ( .A(register__n10372), .Y(register__n10371) );
  BUFx4f_ASAP7_75t_R register___U15014 ( .A(register__n5871), .Y(register__n10372) );
  BUFx4f_ASAP7_75t_R register___U15015 ( .A(register__net117747), .Y(register__net88893) );
  BUFx4f_ASAP7_75t_R register___U15016 ( .A(register__net103649), .Y(register__net88889) );
  BUFx4f_ASAP7_75t_R register___U15017 ( .A(register__net105801), .Y(register__net88885) );
  BUFx6f_ASAP7_75t_R register___U15018 ( .A(register__n10374), .Y(register__n10373) );
  BUFx4f_ASAP7_75t_R register___U15019 ( .A(register__n6879), .Y(register__n10374) );
  BUFx6f_ASAP7_75t_R register___U15020 ( .A(register__n10376), .Y(register__n10375) );
  BUFx4f_ASAP7_75t_R register___U15021 ( .A(register__n8092), .Y(register__n10376) );
  BUFx6f_ASAP7_75t_R register___U15022 ( .A(register__n10378), .Y(register__n10377) );
  BUFx4f_ASAP7_75t_R register___U15023 ( .A(register__n9008), .Y(register__n10378) );
  BUFx6f_ASAP7_75t_R register___U15024 ( .A(register__n10380), .Y(register__n10379) );
  BUFx4f_ASAP7_75t_R register___U15025 ( .A(register__n6116), .Y(register__n10380) );
  BUFx6f_ASAP7_75t_R register___U15026 ( .A(register__n10382), .Y(register__n10381) );
  BUFx4f_ASAP7_75t_R register___U15027 ( .A(register__n7507), .Y(register__n10382) );
  BUFx4f_ASAP7_75t_R register___U15028 ( .A(register__net107984), .Y(register__net88861) );
  BUFx4f_ASAP7_75t_R register___U15029 ( .A(register__net110020), .Y(register__net88857) );
  BUFx6f_ASAP7_75t_R register___U15030 ( .A(register__n10384), .Y(register__n10383) );
  BUFx4f_ASAP7_75t_R register___U15031 ( .A(register__n8137), .Y(register__n10384) );
  BUFx6f_ASAP7_75t_R register___U15032 ( .A(register__n10386), .Y(register__n10385) );
  BUFx4f_ASAP7_75t_R register___U15033 ( .A(register__n8139), .Y(register__n10386) );
  BUFx6f_ASAP7_75t_R register___U15034 ( .A(register__n10388), .Y(register__n10387) );
  BUFx4f_ASAP7_75t_R register___U15035 ( .A(register__n8493), .Y(register__n10388) );
  BUFx6f_ASAP7_75t_R register___U15036 ( .A(register__n10392), .Y(register__n10391) );
  BUFx4f_ASAP7_75t_R register___U15037 ( .A(register__n8151), .Y(register__n10392) );
  BUFx6f_ASAP7_75t_R register___U15038 ( .A(register__n10394), .Y(register__n10393) );
  BUFx4f_ASAP7_75t_R register___U15039 ( .A(register__n7815), .Y(register__n10394) );
  BUFx6f_ASAP7_75t_R register___U15040 ( .A(register__n10396), .Y(register__n10395) );
  BUFx4f_ASAP7_75t_R register___U15041 ( .A(register__n7817), .Y(register__n10396) );
  BUFx6f_ASAP7_75t_R register___U15042 ( .A(register__n10398), .Y(register__n10397) );
  BUFx4f_ASAP7_75t_R register___U15043 ( .A(register__n7529), .Y(register__n10398) );
  BUFx4f_ASAP7_75t_R register___U15044 ( .A(register__net105678), .Y(register__net88821) );
  BUFx4f_ASAP7_75t_R register___U15045 ( .A(register__net103449), .Y(register__net88817) );
  BUFx6f_ASAP7_75t_R register___U15046 ( .A(register__net88814), .Y(register__net88813) );
  BUFx4f_ASAP7_75t_R register___U15047 ( .A(register__net98310), .Y(register__net88814) );
  BUFx6f_ASAP7_75t_R register___U15048 ( .A(register__n10400), .Y(register__n10399) );
  BUFx4f_ASAP7_75t_R register___U15049 ( .A(register__n7225), .Y(register__n10400) );
  BUFx6f_ASAP7_75t_R register___U15050 ( .A(register__n10402), .Y(register__n10401) );
  BUFx4f_ASAP7_75t_R register___U15051 ( .A(register__n7543), .Y(register__n10402) );
  BUFx6f_ASAP7_75t_R register___U15052 ( .A(register__n10404), .Y(register__n10403) );
  BUFx4f_ASAP7_75t_R register___U15053 ( .A(register__n7833), .Y(register__n10404) );
  BUFx6f_ASAP7_75t_R register___U15054 ( .A(register__n10406), .Y(register__n10405) );
  BUFx4f_ASAP7_75t_R register___U15055 ( .A(register__n7234), .Y(register__n10406) );
  BUFx6f_ASAP7_75t_R register___U15056 ( .A(register__n10408), .Y(register__n10407) );
  BUFx4f_ASAP7_75t_R register___U15057 ( .A(register__n7557), .Y(register__n10408) );
  BUFx6f_ASAP7_75t_R register___U15058 ( .A(register__n10410), .Y(register__n10409) );
  BUFx4f_ASAP7_75t_R register___U15059 ( .A(register__n7850), .Y(register__n10410) );
  BUFx6f_ASAP7_75t_R register___U15060 ( .A(register__n10412), .Y(register__n10411) );
  BUFx4f_ASAP7_75t_R register___U15061 ( .A(register__n7857), .Y(register__n10412) );
  BUFx6f_ASAP7_75t_R register___U15062 ( .A(register__n10414), .Y(register__n10413) );
  BUFx4f_ASAP7_75t_R register___U15063 ( .A(register__n7859), .Y(register__n10414) );
  BUFx12f_ASAP7_75t_R register___U15064 ( .A(register__n11891), .Y(register__n11890) );
  BUFx6f_ASAP7_75t_R register___U15065 ( .A(register__n10422), .Y(register__n10421) );
  BUFx4f_ASAP7_75t_R register___U15066 ( .A(register__n6348), .Y(register__n10422) );
  BUFx4f_ASAP7_75t_R register___U15067 ( .A(register__net105782), .Y(register__net88628) );
  BUFx6f_ASAP7_75t_R register___U15068 ( .A(register__n10424), .Y(register__n10423) );
  BUFx4f_ASAP7_75t_R register___U15069 ( .A(register__n9017), .Y(register__n10424) );
  BUFx6f_ASAP7_75t_R register___U15070 ( .A(register__n10427), .Y(register__n10426) );
  BUFx4f_ASAP7_75t_R register___U15071 ( .A(register__n8473), .Y(register__n10427) );
  BUFx6f_ASAP7_75t_R register___U15072 ( .A(register__n10429), .Y(register__n10428) );
  BUFx4f_ASAP7_75t_R register___U15073 ( .A(register__n6926), .Y(register__n10429) );
  BUFx6f_ASAP7_75t_R register___U15074 ( .A(register__n10431), .Y(register__n10430) );
  BUFx4f_ASAP7_75t_R register___U15075 ( .A(register__n6846), .Y(register__n10431) );
  BUFx4f_ASAP7_75t_R register___U15076 ( .A(register__net95340), .Y(register__net88604) );
  BUFx6f_ASAP7_75t_R register___U15077 ( .A(register__n10433), .Y(register__n10432) );
  BUFx4f_ASAP7_75t_R register___U15078 ( .A(register__n6599), .Y(register__n10433) );
  BUFx6f_ASAP7_75t_R register___U15079 ( .A(register__n10437), .Y(register__n10436) );
  BUFx4f_ASAP7_75t_R register___U15080 ( .A(register__n6611), .Y(register__n10437) );
  BUFx4f_ASAP7_75t_R register___U15081 ( .A(register__net105754), .Y(register__net88584) );
  BUFx6f_ASAP7_75t_R register___U15082 ( .A(register__n10441), .Y(register__n10440) );
  BUFx4f_ASAP7_75t_R register___U15083 ( .A(register__n7794), .Y(register__n10441) );
  BUFx6f_ASAP7_75t_R register___U15084 ( .A(register__n10445), .Y(register__n10444) );
  BUFx4f_ASAP7_75t_R register___U15085 ( .A(register__n8859), .Y(register__n10445) );
  BUFx6f_ASAP7_75t_R register___U15086 ( .A(register__n10447), .Y(register__n10446) );
  BUFx4f_ASAP7_75t_R register___U15087 ( .A(register__n8861), .Y(register__n10447) );
  BUFx6f_ASAP7_75t_R register___U15088 ( .A(register__n10449), .Y(register__n10448) );
  BUFx4f_ASAP7_75t_R register___U15089 ( .A(register__n6560), .Y(register__n10449) );
  BUFx6f_ASAP7_75t_R register___U15090 ( .A(register__n10451), .Y(register__n10450) );
  BUFx4f_ASAP7_75t_R register___U15091 ( .A(register__n6332), .Y(register__n10451) );
  BUFx4f_ASAP7_75t_R register___U15092 ( .A(register__net103668), .Y(register__net88548) );
  BUFx6f_ASAP7_75t_R register___U15093 ( .A(register__n10453), .Y(register__n10452) );
  BUFx4f_ASAP7_75t_R register___U15094 ( .A(register__n8068), .Y(register__n10453) );
  BUFx4f_ASAP7_75t_R register___U15095 ( .A(register__n8895), .Y(register__n10455) );
  BUFx6f_ASAP7_75t_R register___U15096 ( .A(register__n10457), .Y(register__n10456) );
  BUFx4f_ASAP7_75t_R register___U15097 ( .A(register__n7473), .Y(register__n10457) );
  BUFx6f_ASAP7_75t_R register___U15098 ( .A(register__n10459), .Y(register__n10458) );
  BUFx4f_ASAP7_75t_R register___U15099 ( .A(register__n7480), .Y(register__n10459) );
  BUFx4f_ASAP7_75t_R register___U15100 ( .A(register__n8953), .Y(register__n10461) );
  BUFx6f_ASAP7_75t_R register___U15101 ( .A(register__n10464), .Y(register__n10463) );
  BUFx4f_ASAP7_75t_R register___U15102 ( .A(register__n7181), .Y(register__n10464) );
  BUFx6f_ASAP7_75t_R register___U15103 ( .A(register__n10466), .Y(register__n10465) );
  BUFx4f_ASAP7_75t_R register___U15104 ( .A(register__n7489), .Y(register__n10466) );
  BUFx6f_ASAP7_75t_R register___U15105 ( .A(register__n10468), .Y(register__n10467) );
  BUFx4f_ASAP7_75t_R register___U15106 ( .A(register__n6378), .Y(register__n10468) );
  BUFx4f_ASAP7_75t_R register___U15107 ( .A(register__net139182), .Y(register__net88504) );
  BUFx4f_ASAP7_75t_R register___U15108 ( .A(register__net101112), .Y(register__net88500) );
  BUFx4f_ASAP7_75t_R register___U15109 ( .A(register__net139166), .Y(register__net88496) );
  BUFx6f_ASAP7_75t_R register___U15110 ( .A(register__n10470), .Y(register__n10469) );
  BUFx4f_ASAP7_75t_R register___U15111 ( .A(register__n3812), .Y(register__n10470) );
  BUFx6f_ASAP7_75t_R register___U15112 ( .A(register__n10472), .Y(register__n10471) );
  BUFx4f_ASAP7_75t_R register___U15113 ( .A(register__n7531), .Y(register__n10472) );
  BUFx6f_ASAP7_75t_R register___U15114 ( .A(register__n10474), .Y(register__n10473) );
  BUFx4f_ASAP7_75t_R register___U15115 ( .A(register__n6657), .Y(register__n10474) );
  BUFx6f_ASAP7_75t_R register___U15116 ( .A(register__n10476), .Y(register__n10475) );
  BUFx4f_ASAP7_75t_R register___U15117 ( .A(register__n8214), .Y(register__n10476) );
  BUFx6f_ASAP7_75t_R register___U15118 ( .A(register__n10478), .Y(register__n10477) );
  BUFx4f_ASAP7_75t_R register___U15119 ( .A(register__n5849), .Y(register__n10478) );
  BUFx4f_ASAP7_75t_R register___U15120 ( .A(register__net106029), .Y(register__net88473) );
  BUFx6f_ASAP7_75t_R register___U15121 ( .A(register__n10480), .Y(register__n10479) );
  BUFx4f_ASAP7_75t_R register___U15122 ( .A(register__n5363), .Y(register__n10480) );
  BUFx6f_ASAP7_75t_R register___U15123 ( .A(register__n10482), .Y(register__n10481) );
  BUFx4f_ASAP7_75t_R register___U15124 ( .A(register__n6072), .Y(register__n10482) );
  BUFx6f_ASAP7_75t_R register___U15125 ( .A(register__n10484), .Y(register__n10483) );
  BUFx4f_ASAP7_75t_R register___U15126 ( .A(register__n5667), .Y(register__n10484) );
  BUFx6f_ASAP7_75t_R register___U15127 ( .A(register__n10486), .Y(register__n10485) );
  BUFx4f_ASAP7_75t_R register___U15128 ( .A(register__n5853), .Y(register__n10486) );
  BUFx6f_ASAP7_75t_R register___U15129 ( .A(register__n10488), .Y(register__n10487) );
  BUFx4f_ASAP7_75t_R register___U15130 ( .A(register__n5859), .Y(register__n10488) );
  BUFx6f_ASAP7_75t_R register___U15131 ( .A(register__n10490), .Y(register__n10489) );
  BUFx4f_ASAP7_75t_R register___U15132 ( .A(register__n7434), .Y(register__n10490) );
  BUFx6f_ASAP7_75t_R register___U15133 ( .A(register__n10492), .Y(register__n10491) );
  BUFx4f_ASAP7_75t_R register___U15134 ( .A(register__n5365), .Y(register__n10492) );
  BUFx6f_ASAP7_75t_R register___U15135 ( .A(register__n10494), .Y(register__n10493) );
  BUFx4f_ASAP7_75t_R register___U15136 ( .A(register__n6862), .Y(register__n10494) );
  BUFx6f_ASAP7_75t_R register___U15137 ( .A(register__n10496), .Y(register__n10495) );
  BUFx4f_ASAP7_75t_R register___U15138 ( .A(register__n8873), .Y(register__n10496) );
  BUFx6f_ASAP7_75t_R register___U15139 ( .A(register__n10498), .Y(register__n10497) );
  BUFx4f_ASAP7_75t_R register___U15140 ( .A(register__n3693), .Y(register__n10498) );
  BUFx4f_ASAP7_75t_R register___U15141 ( .A(register__n8921), .Y(register__n10500) );
  BUFx6f_ASAP7_75t_R register___U15142 ( .A(register__n10504), .Y(register__n10503) );
  BUFx4f_ASAP7_75t_R register___U15143 ( .A(register__n8123), .Y(register__n10504) );
  BUFx4f_ASAP7_75t_R register___U15144 ( .A(register__net98415), .Y(register__net88417) );
  BUFx4f_ASAP7_75t_R register___U15145 ( .A(register__net98396), .Y(register__net88412) );
  BUFx4f_ASAP7_75t_R register___U15146 ( .A(register__n9069), .Y(register__n10506) );
  BUFx4f_ASAP7_75t_R register___U15147 ( .A(register__net114093), .Y(register__net88404) );
  BUFx6f_ASAP7_75t_R register___U15148 ( .A(register__n10508), .Y(register__n10507) );
  BUFx4f_ASAP7_75t_R register___U15149 ( .A(register__n6971), .Y(register__n10508) );
  BUFx6f_ASAP7_75t_R register___U15150 ( .A(register__n10510), .Y(register__n10509) );
  BUFx4f_ASAP7_75t_R register___U15151 ( .A(register__n5855), .Y(register__n10510) );
  BUFx6f_ASAP7_75t_R register___U15152 ( .A(register__n10512), .Y(register__n10511) );
  BUFx4f_ASAP7_75t_R register___U15153 ( .A(register__n6595), .Y(register__n10512) );
  BUFx6f_ASAP7_75t_R register___U15154 ( .A(register__n10514), .Y(register__n10513) );
  BUFx4f_ASAP7_75t_R register___U15155 ( .A(register__n8198), .Y(register__n10514) );
  BUFx6f_ASAP7_75t_R register___U15156 ( .A(register__n10516), .Y(register__n10515) );
  BUFx4f_ASAP7_75t_R register___U15157 ( .A(register__n6603), .Y(register__n10516) );
  BUFx12f_ASAP7_75t_R register___U15158 ( .A(Reg_data[946]), .Y(register__n10519) );
  INVx2_ASAP7_75t_R register___U15159 ( .A(register__n10519), .Y(register__n11845) );
  INVxp67_ASAP7_75t_R register___U15160 ( .A(register__n6284), .Y(register__n11844) );
  INVx1_ASAP7_75t_R register___U15161 ( .A(register__n10363), .Y(register__n10529) );
  AND4x1_ASAP7_75t_R register___U15162 ( .A(register__n7320), .B(register__n7319), .C(register__n3664), .D(register__n2977), .Y(
        n10524) );
  AND4x1_ASAP7_75t_R register___U15163 ( .A(register__n8567), .B(register__n7878), .C(register__n8568), .D(register__n5016), .Y(
        n10522) );
  INVx1_ASAP7_75t_R register___U15164 ( .A(register__n10361), .Y(register__n10554) );
  INVx1_ASAP7_75t_R register___U15165 ( .A(register__n10359), .Y(register__n10574) );
  AND4x1_ASAP7_75t_R register___U15166 ( .A(register__n5701), .B(register__n2158), .C(register__n8572), .D(register__n3988), .Y(
        n10569) );
  AND4x1_ASAP7_75t_R register___U15167 ( .A(register__n6703), .B(register__n8637), .C(register__n6704), .D(register__n4446), .Y(
        n10568) );
  INVx1_ASAP7_75t_R register___U15168 ( .A(register__n10357), .Y(register__n10595) );
  INVx1_ASAP7_75t_R register___U15169 ( .A(register__n9467), .Y(register__n10597) );
  INVx1_ASAP7_75t_R register___U15170 ( .A(register__n10355), .Y(register__n10618) );
  AND4x1_ASAP7_75t_R register___U15171 ( .A(register__n7644), .B(register__n7642), .C(register__n6298), .D(register__n4333), .Y(
        n10612) );
  INVx1_ASAP7_75t_R register___U15172 ( .A(register__n10379), .Y(register__n10639) );
  AND4x1_ASAP7_75t_R register___U15173 ( .A(register__n7005), .B(register__n36), .C(register__n7003), .D(register__n5107), .Y(
        n10633) );
  INVx1_ASAP7_75t_R register___U15174 ( .A(register__n10371), .Y(register__n10661) );
  INVx1_ASAP7_75t_R register___U15175 ( .A(register__n10401), .Y(register__n10682) );
  INVx1_ASAP7_75t_R register___U15176 ( .A(register__n10403), .Y(register__n10684) );
  AND4x1_ASAP7_75t_R register___U15177 ( .A(register__n7603), .B(register__n7602), .C(register__n6299), .D(register__n5798), .Y(
        n10678) );
  INVx1_ASAP7_75t_R register___U15178 ( .A(register__net88821), .Y(register__C6422_net59829) );
  INVx1_ASAP7_75t_R register___U15179 ( .A(register__net88817), .Y(register__C6422_net59833) );
  AND4x1_ASAP7_75t_R register___U15180 ( .A(register__n5376), .B(register__n3996), .C(register__n5378), .D(register__n3017), .Y(
        n10699) );
  AND4x1_ASAP7_75t_R register___U15181 ( .A(register__n9149), .B(register__n9150), .C(register__n8383), .D(register__n5422), .Y(
        n10698) );
  INVx1_ASAP7_75t_R register___U15182 ( .A(register__net88885), .Y(register__C6422_net59855) );
  AND4x1_ASAP7_75t_R register___U15183 ( .A(register__n6194), .B(register__n3910), .C(register__n6196), .D(register__n6195), .Y(
        n10717) );
  INVx1_ASAP7_75t_R register___U15184 ( .A(register__n9553), .Y(register__n10739) );
  INVx1_ASAP7_75t_R register___U15185 ( .A(register__n10409), .Y(register__n10742) );
  AND4x1_ASAP7_75t_R register___U15186 ( .A(register__n4976), .B(register__n705), .C(register__n4975), .D(register__n3530), .Y(
        n10734) );
  INVx1_ASAP7_75t_R register___U15187 ( .A(register__n9505), .Y(register__n10761) );
  INVx1_ASAP7_75t_R register___U15188 ( .A(register__n9507), .Y(register__n10763) );
  INVx1_ASAP7_75t_R register___U15189 ( .A(register__n9509), .Y(register__n10762) );
  INVx1_ASAP7_75t_R register___U15190 ( .A(register__n10373), .Y(register__n10764) );
  INVx1_ASAP7_75t_R register___U15191 ( .A(register__n9527), .Y(register__n10787) );
  INVx1_ASAP7_75t_R register___U15192 ( .A(register__n9557), .Y(register__n10788) );
  AND4x1_ASAP7_75t_R register___U15193 ( .A(register__n7946), .B(register__n4380), .C(register__n3634), .D(register__n7944), .Y(
        n10781) );
  AND4x1_ASAP7_75t_R register___U15194 ( .A(register__n6706), .B(register__n1245), .C(register__n1741), .D(register__n4811), .Y(
        n10780) );
  INVx1_ASAP7_75t_R register___U15195 ( .A(register__net91259), .Y(register__C6422_net59959) );
  INVx1_ASAP7_75t_R register___U15196 ( .A(register__net88857), .Y(register__C6422_net59963) );
  INVx1_ASAP7_75t_R register___U15197 ( .A(register__n10353), .Y(register__n10823) );
  INVx1_ASAP7_75t_R register___U15198 ( .A(register__n9517), .Y(register__n10847) );
  INVx1_ASAP7_75t_R register___U15199 ( .A(register__n10381), .Y(register__n10846) );
  INVx1_ASAP7_75t_R register___U15200 ( .A(register__n10369), .Y(register__n10866) );
  INVx1_ASAP7_75t_R register___U15201 ( .A(register__n9479), .Y(register__n10869) );
  AND4x1_ASAP7_75t_R register___U15202 ( .A(register__n7013), .B(register__n3303), .C(register__n7011), .D(register__n3094), .Y(
        n10861) );
  INVx1_ASAP7_75t_R register___U15203 ( .A(register__n8831), .Y(register__n10893) );
  INVx1_ASAP7_75t_R register___U15204 ( .A(register__n10397), .Y(register__n10892) );
  AND4x1_ASAP7_75t_R register___U15205 ( .A(register__n5229), .B(register__n1858), .C(register__n5228), .D(register__n5230), .Y(
        n10885) );
  AND4x1_ASAP7_75t_R register___U15206 ( .A(register__n8634), .B(register__n8632), .C(register__n8633), .D(register__n4772), .Y(
        n10883) );
  INVx1_ASAP7_75t_R register___U15207 ( .A(register__n10367), .Y(register__n10913) );
  AND4x1_ASAP7_75t_R register___U15208 ( .A(register__n8254), .B(register__n8252), .C(register__n8253), .D(register__n4863), .Y(
        n10906) );
  INVx1_ASAP7_75t_R register___U15209 ( .A(register__n9503), .Y(register__n10933) );
  INVx1_ASAP7_75t_R register___U15210 ( .A(register__n10365), .Y(register__n10955) );
  INVx1_ASAP7_75t_R register___U15211 ( .A(register__n10399), .Y(register__n10979) );
  INVx1_ASAP7_75t_R register___U15212 ( .A(register__n9551), .Y(register__n10981) );
  AND4x1_ASAP7_75t_R register___U15213 ( .A(register__n7313), .B(register__n7312), .C(register__n8381), .D(register__n4344), .Y(
        n10973) );
  INVx1_ASAP7_75t_R register___U15214 ( .A(register__net88913), .Y(register__C6422_net60219) );
  AND4x1_ASAP7_75t_R register___U15215 ( .A(register__n6448), .B(register__n6447), .C(register__n3752), .D(register__n6449), .Y(
        n10996) );
  AND4x1_ASAP7_75t_R register___U15216 ( .A(register__n8628), .B(register__n8627), .C(register__n8626), .D(register__n5061), .Y(
        n10994) );
  INVx1_ASAP7_75t_R register___U15217 ( .A(register__n10405), .Y(register__n11017) );
  INVx1_ASAP7_75t_R register___U15218 ( .A(register__n9565), .Y(register__n11019) );
  INVx1_ASAP7_75t_R register___U15219 ( .A(register__n9537), .Y(register__n11018) );
  INVx1_ASAP7_75t_R register___U15220 ( .A(register__n10411), .Y(register__n11041) );
  INVx1_ASAP7_75t_R register___U15221 ( .A(register__n10391), .Y(register__n11059) );
  AND4x1_ASAP7_75t_R register___U15222 ( .A(register__n7916), .B(register__n7917), .C(register__n7918), .D(register__n4996), .Y(
        n11055) );
  INVx1_ASAP7_75t_R register___U15223 ( .A(register__net88756), .Y(register__C6422_net60324) );
  INVx1_ASAP7_75t_R register___U15224 ( .A(register__net88764), .Y(register__C6422_net60323) );
  INVx1_ASAP7_75t_R register___U15225 ( .A(register__net91255), .Y(register__C6422_net60326) );
  INVx1_ASAP7_75t_R register___U15226 ( .A(register__net88752), .Y(register__C6422_net60328) );
  AND4x1_ASAP7_75t_R register___U15227 ( .A(register__n6428), .B(register__n6429), .C(register__n8035), .D(register__n4712), .Y(
        n11079) );
  INVx1_ASAP7_75t_R register___U15228 ( .A(register__n9539), .Y(register__n11103) );
  INVx1_ASAP7_75t_R register___U15229 ( .A(register__n10389), .Y(register__n11107) );
  AND4x1_ASAP7_75t_R register___U15230 ( .A(register__n6458), .B(register__n6457), .C(register__n6459), .D(register__n2888), .Y(
        n11098) );
  INVx1_ASAP7_75t_R register___U15231 ( .A(register__n9515), .Y(register__n11128) );
  INVx1_ASAP7_75t_R register___U15232 ( .A(register__n10417), .Y(register__n11130) );
  INVx1_ASAP7_75t_R register___U15233 ( .A(register__n10363), .Y(register__n11160) );
  AND4x1_ASAP7_75t_R register___U15234 ( .A(register__n7933), .B(register__n7932), .C(register__n5920), .D(register__n2258), .Y(
        n11156) );
  INVx1_ASAP7_75t_R register___U15235 ( .A(register__n10361), .Y(register__n11179) );
  AND4x1_ASAP7_75t_R register___U15236 ( .A(register__n7883), .B(register__n302), .C(register__n1237), .D(register__n7882), .Y(
        n11174) );
  INVx1_ASAP7_75t_R register___U15237 ( .A(register__n10359), .Y(register__n11201) );
  AND4x1_ASAP7_75t_R register___U15238 ( .A(register__n7926), .B(register__n7927), .C(register__n5694), .D(register__n4683), .Y(
        n11197) );
  AND4x1_ASAP7_75t_R register___U15239 ( .A(register__n7010), .B(register__n7008), .C(register__n7261), .D(register__n4239), .Y(
        n11196) );
  AND4x1_ASAP7_75t_R register___U15240 ( .A(register__n6144), .B(register__n6145), .C(register__n6143), .D(register__n2906), .Y(
        n11195) );
  INVx1_ASAP7_75t_R register___U15241 ( .A(register__n10357), .Y(register__n11225) );
  INVx1_ASAP7_75t_R register___U15242 ( .A(register__n9467), .Y(register__n11226) );
  INVx1_ASAP7_75t_R register___U15243 ( .A(register__n10355), .Y(register__n11245) );
  AND4x1_ASAP7_75t_R register___U15244 ( .A(register__n5923), .B(register__n5921), .C(register__n5518), .D(register__n4436), .Y(
        n11240) );
  INVx1_ASAP7_75t_R register___U15245 ( .A(register__net88889), .Y(register__C6423_net60617) );
  INVx1_ASAP7_75t_R register___U15246 ( .A(register__net88893), .Y(register__C6423_net60643) );
  INVx1_ASAP7_75t_R register___U15247 ( .A(register__net91463), .Y(register__C6423_net60645) );
  AND4x1_ASAP7_75t_R register___U15248 ( .A(register__n7265), .B(register__n1506), .C(register__n7007), .D(register__n4319), .Y(
        n11279) );
  AND4x1_ASAP7_75t_R register___U15249 ( .A(register__n6698), .B(register__n6697), .C(register__n6699), .D(register__n4272), .Y(
        n11278) );
  INVx1_ASAP7_75t_R register___U15250 ( .A(register__n10379), .Y(register__n11304) );
  AND4x1_ASAP7_75t_R register___U15251 ( .A(register__n5925), .B(register__n1508), .C(register__n5924), .D(register__n3919), .Y(
        n11298) );
  AND4x1_ASAP7_75t_R register___U15252 ( .A(register__n6151), .B(register__n6152), .C(register__n6150), .D(register__n2864), .Y(
        n11297) );
  INVx1_ASAP7_75t_R register___U15253 ( .A(register__n10371), .Y(register__n11326) );
  INVx1_ASAP7_75t_R register___U15254 ( .A(register__n10401), .Y(register__n11348) );
  INVx1_ASAP7_75t_R register___U15255 ( .A(register__n10403), .Y(register__n11351) );
  AND4x1_ASAP7_75t_R register___U15256 ( .A(register__n152), .B(register__n6420), .C(register__n1242), .D(register__n4558), .Y(
        n11342) );
  INVx1_ASAP7_75t_R register___U15257 ( .A(register__n9553), .Y(register__n11371) );
  INVx1_ASAP7_75t_R register___U15258 ( .A(register__n10409), .Y(register__n11373) );
  AND4x1_ASAP7_75t_R register___U15259 ( .A(register__n5917), .B(register__n5918), .C(register__n6057), .D(register__n5436), .Y(
        n11366) );
  INVx1_ASAP7_75t_R register___U15260 ( .A(register__n9505), .Y(register__n11392) );
  INVx1_ASAP7_75t_R register___U15261 ( .A(register__n9523), .Y(register__n11391) );
  INVx1_ASAP7_75t_R register___U15262 ( .A(register__n9507), .Y(register__n11394) );
  INVx1_ASAP7_75t_R register___U15263 ( .A(register__n9509), .Y(register__n11393) );
  AND4x1_ASAP7_75t_R register___U15264 ( .A(register__n7301), .B(register__n7302), .C(register__n5842), .D(register__n4700), .Y(
        n11386) );
  INVx1_ASAP7_75t_R register___U15265 ( .A(register__n9541), .Y(register__n11412) );
  INVx1_ASAP7_75t_R register___U15266 ( .A(register__n9557), .Y(register__n11414) );
  AND4x1_ASAP7_75t_R register___U15267 ( .A(register__n6155), .B(register__n6156), .C(register__n5663), .D(register__n5429), .Y(
        n11407) );
  AND4x1_ASAP7_75t_R register___U15268 ( .A(register__n7598), .B(register__n2087), .C(register__n7599), .D(register__n2873), .Y(
        n11406) );
  INVx1_ASAP7_75t_R register___U15269 ( .A(register__n10353), .Y(register__n11434) );
  AND4x1_ASAP7_75t_R register___U15270 ( .A(register__n1482), .B(register__n1610), .C(register__n1369), .D(register__n1061), .Y(
        n11430) );
  INVx1_ASAP7_75t_R register___U15271 ( .A(register__n9517), .Y(register__n11458) );
  INVx1_ASAP7_75t_R register___U15272 ( .A(register__n10381), .Y(register__n11457) );
  INVx1_ASAP7_75t_R register___U15273 ( .A(register__n10369), .Y(register__n11479) );
  INVx1_ASAP7_75t_R register___U15274 ( .A(register__n9479), .Y(register__n11480) );
  AND4x1_ASAP7_75t_R register___U15275 ( .A(register__n6408), .B(register__n6406), .C(register__n7260), .D(register__n4018), .Y(
        n11473) );
  AND4x1_ASAP7_75t_R register___U15276 ( .A(register__n7637), .B(register__n7635), .C(register__n3869), .D(register__n3088), .Y(
        n11472) );
  INVx1_ASAP7_75t_R register___U15277 ( .A(register__n8831), .Y(register__n11504) );
  INVx1_ASAP7_75t_R register___U15278 ( .A(register__n10397), .Y(register__n11502) );
  AND4x1_ASAP7_75t_R register___U15279 ( .A(register__n7270), .B(register__n7269), .C(register__n5519), .D(register__n4704), .Y(
        n11495) );
  AND4x1_ASAP7_75t_R register___U15280 ( .A(register__n5231), .B(register__n5233), .C(register__n2924), .D(register__n4119), .Y(
        n11494) );
  INVx1_ASAP7_75t_R register___U15281 ( .A(register__n10367), .Y(register__n11524) );
  AND4x1_ASAP7_75t_R register___U15282 ( .A(register__n6415), .B(register__n6413), .C(register__n5517), .D(register__n4314), .Y(
        n11518) );
  AND4x1_ASAP7_75t_R register___U15283 ( .A(register__n7880), .B(register__n1464), .C(register__n1504), .D(register__n3054), .Y(
        n11517) );
  AND4x1_ASAP7_75t_R register___U15284 ( .A(register__n7923), .B(register__n7924), .C(register__n6749), .D(register__n784), .Y(
        n11542) );
  INVx1_ASAP7_75t_R register___U15285 ( .A(register__n10365), .Y(register__n11566) );
  AND4x1_ASAP7_75t_R register___U15286 ( .A(register__n8259), .B(register__n8258), .C(register__n7921), .D(register__n4552), .Y(
        n11562) );
  AND4x1_ASAP7_75t_R register___U15287 ( .A(register__n8581), .B(register__n8579), .C(register__n5844), .D(register__n4098), .Y(
        n11561) );
  AND4x1_ASAP7_75t_R register___U15288 ( .A(register__n1341), .B(register__n5696), .C(register__n4640), .D(register__n3202), .Y(
        n11560) );
  INVx1_ASAP7_75t_R register___U15289 ( .A(register__n10399), .Y(register__n11583) );
  INVx1_ASAP7_75t_R register___U15290 ( .A(register__n9551), .Y(register__n11586) );
  INVx1_ASAP7_75t_R register___U15291 ( .A(register__net88861), .Y(register__C6423_net61111) );
  INVx1_ASAP7_75t_R register___U15292 ( .A(register__net91335), .Y(register__C6423_net61113) );
  INVx1_ASAP7_75t_R register___U15293 ( .A(register__net88785), .Y(register__C6423_net61116) );
  INVx1_ASAP7_75t_R register___U15294 ( .A(register__net91331), .Y(register__C6423_net61115) );
  AND4x1_ASAP7_75t_R register___U15295 ( .A(register__n1407), .B(register__n6159), .C(register__n1874), .D(register__n4562), .Y(
        n11601) );
  AND4x1_ASAP7_75t_R register___U15296 ( .A(register__n7876), .B(register__n1168), .C(register__n7877), .D(register__n3591), .Y(
        n11600) );
  INVx1_ASAP7_75t_R register___U15297 ( .A(register__n10405), .Y(register__n11622) );
  INVx1_ASAP7_75t_R register___U15298 ( .A(register__n9565), .Y(register__n11625) );
  INVx1_ASAP7_75t_R register___U15299 ( .A(register__n9537), .Y(register__n11624) );
  INVx1_ASAP7_75t_R register___U15300 ( .A(register__n10411), .Y(register__n11643) );
  AND4x1_ASAP7_75t_R register___U15301 ( .A(register__n1083), .B(register__n7653), .C(register__n3466), .D(register__n3111), .Y(
        n11638) );
  INVx1_ASAP7_75t_R register___U15302 ( .A(register__n10391), .Y(register__n11663) );
  INVx1_ASAP7_75t_R register___U15303 ( .A(register__n10419), .Y(register__n11665) );
  INVx1_ASAP7_75t_R register___U15304 ( .A(register__n9539), .Y(register__n11685) );
  AND4x1_ASAP7_75t_R register___U15305 ( .A(register__n6708), .B(register__n6709), .C(register__n6058), .D(register__n5605), .Y(
        n11679) );
  INVx1_ASAP7_75t_R register___U15306 ( .A(register__n7846), .Y(register__n11706) );
  INVx1_ASAP7_75t_R register___U15307 ( .A(register__n10415), .Y(register__n11705) );
  INVx1_ASAP7_75t_R register___U15308 ( .A(register__n9515), .Y(register__n11707) );
  AND4x1_ASAP7_75t_R register___U15309 ( .A(register__n7056), .B(register__n7058), .C(register__n1761), .D(register__n4171), .Y(
        n11700) );
  INVx3_ASAP7_75t_R register___U15310 ( .A(register__n12185), .Y(register__n12173) );
  INVx3_ASAP7_75t_R register___U15311 ( .A(register__net63038), .Y(register__net63004) );
  INVx3_ASAP7_75t_R register___U15312 ( .A(register__net63032), .Y(register__net62988) );
  INVx3_ASAP7_75t_R register___U15313 ( .A(register__net64028), .Y(register__net63998) );
  INVx3_ASAP7_75t_R register___U15314 ( .A(register__net63024), .Y(register__net62992) );
  INVx3_ASAP7_75t_R register___U15315 ( .A(register__net63024), .Y(register__net62986) );
  INVx3_ASAP7_75t_R register___U15316 ( .A(register__n12297), .Y(register__n12283) );
  INVx3_ASAP7_75t_R register___U15317 ( .A(register__n12295), .Y(register__n12280) );
  INVx3_ASAP7_75t_R register___U15318 ( .A(register__n12307), .Y(register__n12292) );
  INVx3_ASAP7_75t_R register___U15319 ( .A(register__net62870), .Y(register__net62836) );
  BUFx12f_ASAP7_75t_R register___U15320 ( .A(register__n5530), .Y(register__n11758) );
  AO22x1_ASAP7_75t_R register___U15321 ( .A1(register__n12387), .A2(register__n1418), .B1(register__n11844), .B2(register__n1414), 
        .Y(register__n12988) );
  INVx3_ASAP7_75t_R register___U15322 ( .A(register__n12381), .Y(register__n12367) );
  INVx2_ASAP7_75t_R register___U15323 ( .A(register__net64056), .Y(register__net64002) );
  INVx3_ASAP7_75t_R register___U15324 ( .A(register__net64724), .Y(register__net64670) );
  INVx2_ASAP7_75t_R register___U15325 ( .A(register__n12140), .Y(register__n12123) );
  INVx3_ASAP7_75t_R register___U15326 ( .A(register__n12139), .Y(register__n12122) );
  INVx3_ASAP7_75t_R register___U15327 ( .A(register__net63026), .Y(register__net62994) );
  INVx2_ASAP7_75t_R register___U15328 ( .A(register__net64706), .Y(register__net64674) );
  INVx3_ASAP7_75t_R register___U15329 ( .A(register__n12045), .Y(register__n12031) );
  INVx3_ASAP7_75t_R register___U15330 ( .A(register__n12011), .Y(register__n11994) );
  INVx3_ASAP7_75t_R register___U15331 ( .A(register__n12275), .Y(register__n12261) );
  INVx3_ASAP7_75t_R register___U15332 ( .A(register__n12042), .Y(register__n12026) );
  INVx2_ASAP7_75t_R register___U15333 ( .A(register__n12010), .Y(register__n11993) );
  INVx3_ASAP7_75t_R register___U15334 ( .A(register__n12004), .Y(register__n11988) );
  INVx2_ASAP7_75t_R register___U15335 ( .A(register__n12047), .Y(register__n12030) );
  INVx2_ASAP7_75t_R register___U15336 ( .A(register__n12039), .Y(register__n12024) );
  INVx3_ASAP7_75t_R register___U15337 ( .A(register__n12036), .Y(register__n12021) );
  INVx3_ASAP7_75t_R register___U15338 ( .A(register__n12038), .Y(register__n12023) );
  INVx3_ASAP7_75t_R register___U15339 ( .A(register__n12324), .Y(register__n12310) );
  INVx2_ASAP7_75t_R register___U15340 ( .A(register__n12046), .Y(register__n12029) );
  INVx2_ASAP7_75t_R register___U15341 ( .A(register__n12441), .Y(register__n12425) );
  INVx3_ASAP7_75t_R register___U15342 ( .A(register__n12437), .Y(register__n12420) );
  INVx3_ASAP7_75t_R register___U15343 ( .A(register__net63036), .Y(register__net63002) );
  BUFx6f_ASAP7_75t_R register___U15344 ( .A(register__net122406), .Y(register__net63288) );
  BUFx12f_ASAP7_75t_R register___U15345 ( .A(register__net103248), .Y(register__net63300) );
  INVx3_ASAP7_75t_R register___U15346 ( .A(register__net63288), .Y(register__net63254) );
  BUFx6f_ASAP7_75t_R register___U15347 ( .A(register__net92027), .Y(register__net63272) );
  INVx3_ASAP7_75t_R register___U15348 ( .A(register__net64892), .Y(register__net64856) );
  BUFx12f_ASAP7_75t_R register___U15349 ( .A(register__net62884), .Y(register__net62848) );
  BUFx6f_ASAP7_75t_R register___U15350 ( .A(register__n12108), .Y(register__n12100) );
  INVx3_ASAP7_75t_R register___U15351 ( .A(register__n12014), .Y(register__n11996) );
  BUFx12f_ASAP7_75t_R register___U15352 ( .A(register__n3596), .Y(register__n12334) );
  INVx3_ASAP7_75t_R register___U15353 ( .A(register__n12013), .Y(register__n11995) );
  BUFx6f_ASAP7_75t_R register___U15354 ( .A(register__net100610), .Y(register__net63380) );
  BUFx6f_ASAP7_75t_R register___U15355 ( .A(register__net133741), .Y(register__net64386) );
  INVx2_ASAP7_75t_R register___U15356 ( .A(register__n12009), .Y(register__n11992) );
  BUFx12f_ASAP7_75t_R register___U15357 ( .A(register__n12449), .Y(register__n12448) );
  INVx3_ASAP7_75t_R register___U15358 ( .A(register__net62868), .Y(register__net62834) );
  INVx3_ASAP7_75t_R register___U15359 ( .A(register__net64800), .Y(register__net64766) );
  BUFx6f_ASAP7_75t_R register___U15360 ( .A(register__n4595), .Y(register__n12043) );
  BUFx12f_ASAP7_75t_R register___U15361 ( .A(register__n4865), .Y(register__n12048) );
  INVx3_ASAP7_75t_R register___U15362 ( .A(register__n12043), .Y(register__n12027) );
  BUFx6f_ASAP7_75t_R register___U15363 ( .A(register__n5223), .Y(register__n12474) );
  INVx3_ASAP7_75t_R register___U15364 ( .A(register__n12474), .Y(register__n12459) );
  BUFx12f_ASAP7_75t_R register___U15365 ( .A(register__n3650), .Y(register__n12154) );
  BUFx12f_ASAP7_75t_R register___U15366 ( .A(register__n3188), .Y(register__n11965) );
  BUFx12f_ASAP7_75t_R register___U15367 ( .A(register__n3537), .Y(register__n12481) );
  BUFx12f_ASAP7_75t_R register___U15368 ( .A(register__n3845), .Y(register__n12189) );
  OR5x1_ASAP7_75t_R register___U15369 ( .A(register__n430), .B(register__n2222), .C(register__n5441), .D(register__n244), .E(register__n821), .Y(register__n12508) );
  INVx1_ASAP7_75t_R register___U15370 ( .A(rst), .Y(register__n12516) );
  OR2x2_ASAP7_75t_R register___U15371 ( .A(register__n6724), .B(register__n1507), .Y(register__net61445) );


    NOR3x1_ASAP7_75t_R imm_gen___U2 ( .A(inst[6]), .B(imm_gen__n24), .C(imm_gen__n98), .Y(imm_gen__n4) );
  INVx2_ASAP7_75t_R imm_gen___U3 ( .A(imm_gen__n80), .Y(imm_gen__n115) );
  BUFx6f_ASAP7_75t_R imm_gen___U4 ( .A(imm_gen__n11), .Y(imm_gen__n75) );
  NAND2xp33_ASAP7_75t_R imm_gen___U5 ( .A(imm_gen__n11), .B(imm_gen__n17), .Y(imm_gen__n7) );
  BUFx12f_ASAP7_75t_R imm_gen___U6 ( .A(imm_gen__n75), .Y(imm_gen__n74) );
  NAND2x1p5_ASAP7_75t_R imm_gen___U7 ( .A(inst[5]), .B(imm_gen__imm_gen__n102), .Y(imm_gen__n1) );
  NAND2xp5_ASAP7_75t_R imm_gen___U8 ( .A(imm_gen__n72), .B(imm_gen__n2), .Y(imm_gen__n14) );
  INVx1_ASAP7_75t_R imm_gen___U9 ( .A(imm_gen__n1), .Y(imm_gen__n2) );
  INVx3_ASAP7_75t_R imm_gen___U10 ( .A(imm_gen__n111), .Y(imm_gen__n43) );
  INVx2_ASAP7_75t_R imm_gen___U11 ( .A(inst[4]), .Y(imm_gen__n102) );
  INVx3_ASAP7_75t_R imm_gen___U12 ( .A(imm_gen__n24), .Y(imm_gen__n72) );
  INVx3_ASAP7_75t_R imm_gen___U13 ( .A(imm_gen__n43), .Y(imm_gen__n82) );
  NAND2xp33_ASAP7_75t_R imm_gen___U14 ( .A(imm_gen__n11), .B(imm_gen__n17), .Y(imm_gen__n10) );
  NAND2x2_ASAP7_75t_R imm_gen___U15 ( .A(imm_gen__imm_gen__n110), .B(imm_gen__n68), .Y(imm_gen__n11) );
  NAND2xp5_ASAP7_75t_R imm_gen___U16 ( .A(inst[22]), .B(imm_gen__n10), .Y(imm_gen__n3) );
  INVx2_ASAP7_75t_R imm_gen___U17 ( .A(imm_gen__n50), .Y(imm[2]) );
  NAND2x2_ASAP7_75t_R imm_gen___U18 ( .A(imm_gen__n16), .B(imm_gen__n4), .Y(imm_gen__n17) );
  INVx6_ASAP7_75t_R imm_gen___U19 ( .A(imm_gen__n84), .Y(imm_gen__n16) );
  OA211x2_ASAP7_75t_R imm_gen___U20 ( .A1(imm_gen__n120), .A2(imm_gen__n80), .B(inst[31]), .C(imm_gen__n68), .Y(imm_gen__n5)
         );
  OR3x1_ASAP7_75t_R imm_gen___U21 ( .A(inst[6]), .B(imm_gen__n24), .C(imm_gen__n98), .Y(imm_gen__n20) );
  CKINVDCx10_ASAP7_75t_R imm_gen___U22 ( .A(imm_gen__n67), .Y(imm_gen__n84) );
  BUFx12f_ASAP7_75t_R imm_gen___U23 ( .A(imm_gen__n68), .Y(imm_gen__n67) );
  NOR2x1p5_ASAP7_75t_R imm_gen___U24 ( .A(imm_gen__n84), .B(imm_gen__n83), .Y(imm_gen__n111) );
  NOR2x2_ASAP7_75t_R imm_gen___U25 ( .A(imm_gen__n80), .B(imm_gen__n23), .Y(imm_gen__n83) );
  BUFx6f_ASAP7_75t_R imm_gen___U26 ( .A(imm_gen__n117), .Y(imm_gen__n41) );
  AND2x2_ASAP7_75t_R imm_gen___U27 ( .A(imm_gen__n13), .B(imm_gen__n20), .Y(imm_gen__n119) );
  INVxp33_ASAP7_75t_R imm_gen___U28 ( .A(imm_gen__n20), .Y(imm_gen__n99) );
  INVxp67_ASAP7_75t_R imm_gen___U29 ( .A(imm_gen__n42), .Y(imm[3]) );
  HB1xp67_ASAP7_75t_R imm_gen___U30 ( .A(imm_gen__n139), .Y(imm_gen__n42) );
  NOR2xp33_ASAP7_75t_R imm_gen___U31 ( .A(inst[6]), .B(imm_gen__n14), .Y(imm_gen__n6) );
  NAND2xp33_ASAP7_75t_R imm_gen___U32 ( .A(imm_gen__n11), .B(imm_gen__n17), .Y(imm_gen__n8) );
  INVx1_ASAP7_75t_R imm_gen___U33 ( .A(imm_gen__n132), .Y(imm[11]) );
  INVx6_ASAP7_75t_R imm_gen___U34 ( .A(imm_gen__n65), .Y(imm_gen__n80) );
  BUFx3_ASAP7_75t_R imm_gen___U35 ( .A(imm_gen__n118), .Y(imm_gen__n40) );
  INVxp67_ASAP7_75t_R imm_gen___U36 ( .A(imm_gen__n110), .Y(imm_gen__n56) );
  INVx3_ASAP7_75t_R imm_gen___U37 ( .A(imm_gen__n21), .Y(imm_gen__n23) );
  AND2x4_ASAP7_75t_R imm_gen___U38 ( .A(inst[0]), .B(inst[1]), .Y(imm_gen__n117) );
  INVxp67_ASAP7_75t_R imm_gen___U39 ( .A(imm_gen__n45), .Y(imm_gen__n22) );
  OR2x2_ASAP7_75t_R imm_gen___U40 ( .A(imm_gen__n26), .B(imm_gen__n43), .Y(imm_gen__n12) );
  OR2x2_ASAP7_75t_R imm_gen___U41 ( .A(imm_gen__n26), .B(imm_gen__n43), .Y(imm_gen__n15) );
  INVx2_ASAP7_75t_R imm_gen___U42 ( .A(imm_gen__n43), .Y(imm_gen__n44) );
  INVxp67_ASAP7_75t_R imm_gen___U43 ( .A(imm_gen__n12), .Y(imm[20]) );
  INVxp67_ASAP7_75t_R imm_gen___U44 ( .A(imm_gen__n12), .Y(imm[21]) );
  INVxp67_ASAP7_75t_R imm_gen___U45 ( .A(imm_gen__n15), .Y(imm[31]) );
  INVxp67_ASAP7_75t_R imm_gen___U46 ( .A(imm_gen__n15), .Y(imm[22]) );
  INVxp67_ASAP7_75t_R imm_gen___U47 ( .A(imm_gen__n15), .Y(imm[23]) );
  INVxp67_ASAP7_75t_R imm_gen___U48 ( .A(imm_gen__n15), .Y(imm[24]) );
  INVxp67_ASAP7_75t_R imm_gen___U49 ( .A(imm_gen__n15), .Y(imm[27]) );
  INVxp67_ASAP7_75t_R imm_gen___U50 ( .A(imm_gen__n15), .Y(imm[25]) );
  INVxp67_ASAP7_75t_R imm_gen___U51 ( .A(imm_gen__n15), .Y(imm[26]) );
  INVxp67_ASAP7_75t_R imm_gen___U52 ( .A(imm_gen__n15), .Y(imm[28]) );
  INVxp67_ASAP7_75t_R imm_gen___U53 ( .A(imm_gen__n12), .Y(imm[29]) );
  HB1xp67_ASAP7_75t_R imm_gen___U54 ( .A(imm_gen__n33), .Y(imm[18]) );
  INVx1_ASAP7_75t_R imm_gen___U55 ( .A(imm_gen__n76), .Y(imm[30]) );
  INVx2_ASAP7_75t_R imm_gen___U56 ( .A(imm_gen__n122), .Y(imm_gen__n76) );
  INVx3_ASAP7_75t_R imm_gen___U57 ( .A(imm_gen__n12), .Y(imm_gen__imm_gen__n122) );
  OR2x2_ASAP7_75t_R imm_gen___U58 ( .A(inst[6]), .B(imm_gen__n14), .Y(imm_gen__n13) );
  INVx1_ASAP7_75t_R imm_gen___U59 ( .A(imm_gen__n103), .Y(imm_gen__n18) );
  AOI21x1_ASAP7_75t_R imm_gen___U60 ( .A1(imm_gen__n47), .A2(inst[11]), .B(imm_gen__n108), .Y(imm_gen__n138) );
  INVx1_ASAP7_75t_R imm_gen___U61 ( .A(imm_gen__n106), .Y(imm_gen__n19) );
  BUFx3_ASAP7_75t_R imm_gen___U62 ( .A(imm_gen__n140), .Y(imm_gen__n50) );
  CKINVDCx10_ASAP7_75t_R imm_gen___U63 ( .A(imm_gen__n74), .Y(imm_gen__n85) );
  HB1xp67_ASAP7_75t_R imm_gen___U64 ( .A(imm_gen__n30), .Y(imm_gen__n33) );
  BUFx3_ASAP7_75t_R imm_gen___U65 ( .A(imm_gen__n138), .Y(imm_gen__n39) );
  NOR2xp33_ASAP7_75t_R imm_gen___U66 ( .A(imm_gen__n25), .B(imm_gen__n43), .Y(imm_gen__n134) );
  HB1xp67_ASAP7_75t_R imm_gen___U67 ( .A(imm_gen__n13), .Y(imm_gen__n101) );
  AND2x2_ASAP7_75t_R imm_gen___U68 ( .A(imm_gen__n56), .B(imm_gen__n22), .Y(imm_gen__n21) );
  BUFx6f_ASAP7_75t_R imm_gen___U69 ( .A(imm_gen__n119), .Y(imm_gen__n66) );
  BUFx12f_ASAP7_75t_R imm_gen___U70 ( .A(imm_gen__n66), .Y(imm_gen__n65) );
  INVx4_ASAP7_75t_R imm_gen___U71 ( .A(imm_gen__n45), .Y(imm_gen__n79) );
  HB1xp67_ASAP7_75t_R imm_gen___U72 ( .A(imm_gen__n31), .Y(imm_gen__n30) );
  HB1xp67_ASAP7_75t_R imm_gen___U73 ( .A(imm_gen__n125), .Y(imm_gen__n31) );
  OR2x2_ASAP7_75t_R imm_gen___U74 ( .A(n2), .B(inst[2]), .Y(imm_gen__n24) );
  INVxp33_ASAP7_75t_R imm_gen___U75 ( .A(n2), .Y(imm_gen__n97) );
  CKINVDCx20_ASAP7_75t_R imm_gen___U76 ( .A(inst[29]), .Y(imm_gen__n25) );
  HB1xp67_ASAP7_75t_R imm_gen___U77 ( .A(imm_gen__n137), .Y(imm[5]) );
  CKINVDCx20_ASAP7_75t_R imm_gen___U78 ( .A(inst[31]), .Y(imm_gen__n26) );
  HB1xp67_ASAP7_75t_R imm_gen___U79 ( .A(inst[2]), .Y(imm_gen__n27) );
  INVxp33_ASAP7_75t_R imm_gen___U80 ( .A(imm_gen__n97), .Y(imm_gen__n28) );
  AND3x1_ASAP7_75t_R imm_gen___U81 ( .A(inst[5]), .B(imm_gen__n102), .C(imm_gen__n72), .Y(imm_gen__n29) );
  AND2x2_ASAP7_75t_R imm_gen___U82 ( .A(inst[6]), .B(imm_gen__n29), .Y(imm_gen__n113) );
  AO21x1_ASAP7_75t_R imm_gen___U83 ( .A1(inst[18]), .A2(imm_gen__n85), .B(imm_gen__n121), .Y(imm_gen__n125) );
  BUFx2_ASAP7_75t_R imm_gen___U84 ( .A(imm_gen__n124), .Y(imm[19]) );
  AO21x1_ASAP7_75t_R imm_gen___U85 ( .A1(inst[19]), .A2(imm_gen__n85), .B(imm_gen__n121), .Y(imm_gen__n124) );
  BUFx2_ASAP7_75t_R imm_gen___U86 ( .A(imm_gen__n126), .Y(imm[17]) );
  AO21x1_ASAP7_75t_R imm_gen___U87 ( .A1(inst[17]), .A2(imm_gen__n85), .B(imm_gen__n5), .Y(imm_gen__n126) );
  BUFx2_ASAP7_75t_R imm_gen___U88 ( .A(imm_gen__n127), .Y(imm[16]) );
  AO21x1_ASAP7_75t_R imm_gen___U89 ( .A1(inst[16]), .A2(imm_gen__n85), .B(imm_gen__n5), .Y(imm_gen__n127) );
  BUFx2_ASAP7_75t_R imm_gen___U90 ( .A(imm_gen__n133), .Y(imm[10]) );
  BUFx2_ASAP7_75t_R imm_gen___U91 ( .A(imm_gen__n129), .Y(imm[14]) );
  AO21x1_ASAP7_75t_R imm_gen___U92 ( .A1(inst[14]), .A2(imm_gen__n85), .B(imm_gen__n121), .Y(imm_gen__n129) );
  INVx6_ASAP7_75t_R imm_gen___U93 ( .A(imm_gen__n47), .Y(imm_gen__n81) );
  BUFx12f_ASAP7_75t_R imm_gen___U94 ( .A(imm_gen__n113), .Y(imm_gen__n45) );
  BUFx2_ASAP7_75t_R imm_gen___U95 ( .A(imm_gen__n114), .Y(imm_gen__n46) );
  BUFx6f_ASAP7_75t_R imm_gen___U96 ( .A(inst[7]), .Y(imm_gen__n112) );
  BUFx12f_ASAP7_75t_R imm_gen___U97 ( .A(imm_gen__n48), .Y(imm_gen__n47) );
  BUFx12f_ASAP7_75t_R imm_gen___U98 ( .A(imm_gen__n109), .Y(imm_gen__n48) );
  BUFx2_ASAP7_75t_R imm_gen___U99 ( .A(imm_gen__n6), .Y(imm_gen__n49) );
  BUFx2_ASAP7_75t_R imm_gen___U100 ( .A(imm_gen__n134), .Y(imm[9]) );
  BUFx2_ASAP7_75t_R imm_gen___U101 ( .A(imm_gen__n100), .Y(imm_gen__n52) );
  BUFx2_ASAP7_75t_R imm_gen___U102 ( .A(imm_gen__n58), .Y(imm_gen__n53) );
  BUFx4f_ASAP7_75t_R imm_gen___U103 ( .A(imm_gen__n59), .Y(imm[0]) );
  BUFx3_ASAP7_75t_R imm_gen___U104 ( .A(imm_gen__n60), .Y(imm_gen__n59) );
  BUFx2_ASAP7_75t_R imm_gen___U105 ( .A(imm_gen__n128), .Y(imm[15]) );
  AO21x1_ASAP7_75t_R imm_gen___U106 ( .A1(inst[15]), .A2(imm_gen__n85), .B(imm_gen__n5), .Y(imm_gen__n128) );
  AND5x1_ASAP7_75t_R imm_gen___U107 ( .A(inst[6]), .B(inst[5]), .C(imm_gen__n28), .D(imm_gen__n27), .E(
        n102), .Y(imm_gen__n110) );
  AND2x2_ASAP7_75t_R imm_gen___U108 ( .A(inst[24]), .B(imm_gen__n8), .Y(imm_gen__n108) );
  INVx1_ASAP7_75t_R imm_gen___U109 ( .A(imm_gen__n39), .Y(imm[4]) );
  AND2x2_ASAP7_75t_R imm_gen___U110 ( .A(imm_gen__n99), .B(inst[20]), .Y(imm_gen__n100) );
  INVx1_ASAP7_75t_R imm_gen___U111 ( .A(imm_gen__n52), .Y(imm_gen__n58) );
  BUFx2_ASAP7_75t_R imm_gen___U112 ( .A(imm_gen__n142), .Y(imm_gen__n60) );
  BUFx2_ASAP7_75t_R imm_gen___U113 ( .A(imm_gen__n130), .Y(imm[13]) );
  AO21x1_ASAP7_75t_R imm_gen___U114 ( .A1(inst[13]), .A2(imm_gen__n85), .B(imm_gen__n121), .Y(imm_gen__n130) );
  AND2x2_ASAP7_75t_R imm_gen___U115 ( .A(inst[23]), .B(imm_gen__n7), .Y(imm_gen__n106) );
  OA21x2_ASAP7_75t_R imm_gen___U116 ( .A1(imm_gen__n81), .A2(imm_gen__n107), .B(imm_gen__n19), .Y(imm_gen__n139) );
  INVx1_ASAP7_75t_R imm_gen___U117 ( .A(imm_gen__n112), .Y(imm_gen__n63) );
  INVx1_ASAP7_75t_R imm_gen___U118 ( .A(imm_gen__n112), .Y(imm_gen__n64) );
  BUFx12f_ASAP7_75t_R imm_gen___U119 ( .A(imm_gen__n41), .Y(imm_gen__n68) );
  BUFx2_ASAP7_75t_R imm_gen___U120 ( .A(imm_gen__n135), .Y(imm[7]) );
  OA21x2_ASAP7_75t_R imm_gen___U121 ( .A1(imm_gen__n81), .A2(imm_gen__n105), .B(imm_gen__n3), .Y(imm_gen__n140) );
  OA22x2_ASAP7_75t_R imm_gen___U122 ( .A1(imm_gen__n84), .A2(imm_gen__n40), .B1(imm_gen__n11), .B2(imm_gen__imm_gen__n116), .Y(imm_gen__n132)
         );
  INVx1_ASAP7_75t_R imm_gen___U123 ( .A(inst[20]), .Y(imm_gen__n116) );
  BUFx2_ASAP7_75t_R imm_gen___U124 ( .A(imm_gen__n136), .Y(imm[6]) );
  INVx2_ASAP7_75t_R imm_gen___U125 ( .A(imm_gen__n79), .Y(imm_gen__n120) );
  BUFx6f_ASAP7_75t_R imm_gen___U126 ( .A(inst[5]), .Y(imm_gen__n98) );
  BUFx2_ASAP7_75t_R imm_gen___U127 ( .A(imm_gen__n131), .Y(imm[12]) );
  AO21x1_ASAP7_75t_R imm_gen___U128 ( .A1(inst[12]), .A2(imm_gen__n85), .B(imm_gen__n5), .Y(imm_gen__n131) );
  AND2x2_ASAP7_75t_R imm_gen___U129 ( .A(inst[21]), .B(imm_gen__n7), .Y(imm_gen__n103) );
  OA21x2_ASAP7_75t_R imm_gen___U130 ( .A1(imm_gen__n81), .A2(imm_gen__n104), .B(imm_gen__n18), .Y(imm_gen__n141) );
  INVx1_ASAP7_75t_R imm_gen___U131 ( .A(imm_gen__n141), .Y(imm[1]) );
  OA21x2_ASAP7_75t_R imm_gen___U132 ( .A1(imm_gen__n120), .A2(imm_gen__n49), .B(imm_gen__n41), .Y(imm_gen__n109) );
  OA211x2_ASAP7_75t_R imm_gen___U133 ( .A1(imm_gen__n120), .A2(imm_gen__n80), .B(inst[31]), .C(imm_gen__n68), .Y(
        n121) );
  O2A1O1Ixp33_ASAP7_75t_R imm_gen___U134 ( .A1(imm_gen__n64), .A2(imm_gen__n101), .B(imm_gen__n53), .C(imm_gen__n84), .Y(
        n142) );
  INVx1_ASAP7_75t_R imm_gen___U135 ( .A(inst[8]), .Y(imm_gen__n104) );
  INVx1_ASAP7_75t_R imm_gen___U136 ( .A(inst[9]), .Y(imm_gen__n105) );
  INVx1_ASAP7_75t_R imm_gen___U137 ( .A(inst[10]), .Y(imm_gen__n107) );
  AND2x2_ASAP7_75t_R imm_gen___U138 ( .A(inst[25]), .B(imm_gen__n44), .Y(imm_gen__n137) );
  AND2x2_ASAP7_75t_R imm_gen___U139 ( .A(inst[26]), .B(imm_gen__n82), .Y(imm_gen__n136) );
  AND2x2_ASAP7_75t_R imm_gen___U140 ( .A(inst[27]), .B(imm_gen__n82), .Y(imm_gen__n135) );
  AND2x2_ASAP7_75t_R imm_gen___U141 ( .A(inst[28]), .B(imm_gen__n82), .Y(imm[8]) );
  AND2x2_ASAP7_75t_R imm_gen___U142 ( .A(inst[30]), .B(imm_gen__n44), .Y(imm_gen__n133) );
  INVx1_ASAP7_75t_R imm_gen___U143 ( .A(inst[31]), .Y(imm_gen__n114) );
  OA22x2_ASAP7_75t_R imm_gen___U144 ( .A1(imm_gen__n115), .A2(imm_gen__n46), .B1(imm_gen__n79), .B2(imm_gen__n63), .Y(imm_gen__n118)
         );



  BUFx4f_ASAP7_75t_R ID___U1 ( .A(n65), .Y(ID__n4) );
  INVx4_ASAP7_75t_R ID___U2 ( .A(ID__n6), .Y(ID__n5) );
  INVx2_ASAP7_75t_R ID___U3 ( .A(WB_write_back_data[3]), .Y(ID__n6) );
  INVxp67_ASAP7_75t_R ID___U4 ( .A(IF_ID_inst[3]), .Y(ID__n1) );
  INVx1_ASAP7_75t_R ID___U5 ( .A(ID__n10), .Y(ID__n9) );
  INVx1_ASAP7_75t_R ID___U6 ( .A(n109), .Y(ID__n10) );
  INVx4_ASAP7_75t_R ID___U7 ( .A(n64), .Y(ID__n12) );
  BUFx4f_ASAP7_75t_R ID___U8 ( .A(WB_write_back_data[18]), .Y(ID__n3) );
  INVx1_ASAP7_75t_R ID___U9 ( .A(ID__n1), .Y(ID__n2) );
  INVx6_ASAP7_75t_R ID___U10 ( .A(ID__n12), .Y(ID__n11) );
  CKINVDCx10_ASAP7_75t_R ID___U11 ( .A(ID__n8), .Y(ID__n7) );
  CKINVDCx10_ASAP7_75t_R ID___U12 ( .A(WB_write_back_data[4]), .Y(ID__n8) );

  DFFASRHQNx1_ASAP7_75t_R ID_EX___ALUSrc_out_reg ( .D(ID_EX__n177), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n738) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___RegWrite_out_reg ( .D(ID_EX__n5), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__ID_EX__n569), .QN(ID_EX__n739) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_25_ ( .D(ID_EX__n14), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n778) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_22_ ( .D(ID_EX__n46), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n781) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_21_ ( .D(ID_EX__n33), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n782) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_20_ ( .D(ID_EX__n45), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n783) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_18_ ( .D(ID_EX__n43), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n785) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_16_ ( .D(ID_EX__n41), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n787) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_8_ ( .D(ID_EX__n64), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n795) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_6_ ( .D(ID_EX__n68), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n797) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_5_ ( .D(ID_EX__n76), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n798) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_4_ ( .D(ID_EX__n32), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n799) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_3_ ( .D(ID_EX__n48), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n800) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_2_ ( .D(ID_EX__n71), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n801) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_1_ ( .D(ID_EX__n38), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n802) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_0_ ( .D(ID_EX__n67), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n803) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_31_ ( .D(ID_EX__n131), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n804) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_30_ ( .D(ID_EX__n17), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n805) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_29_ ( .D(ID_EX__n145), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n806) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_28_ ( .D(ID_EX__n150), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[28]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_27_ ( .D(ID_EX__n211), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[27]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_26_ ( .D(ID_EX__n154), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[26]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_25_ ( .D(ID_EX__n174), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[25]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_24_ ( .D(ID_EX__n133), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[24]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_23_ ( .D(ID_EX__n134), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[23]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_22_ ( .D(ID_EX__n135), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[22]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_21_ ( .D(ID_EX__n137), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[21]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_20_ ( .D(ID_EX__n142), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[20]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_19_ ( .D(ID_EX__n143), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n807) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_18_ ( .D(ID_EX__n24), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[18]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_17_ ( .D(ID_EX__n146), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[17]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_16_ ( .D(ID_EX__n151), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[16]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_15_ ( .D(ID_EX__n175), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n808) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_14_ ( .D(ID_EX__n155), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[14]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_13_ ( .D(ID_EX__n185), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[13]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_12_ ( .D(ID_EX__n285), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[12]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_11_ ( .D(ID_EX__n218), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n809) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_10_ ( .D(ID_EX__n13), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[10]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_9_ ( .D(ID_EX__n171), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[9]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_8_ ( .D(ID_EX__n258), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[8]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_7_ ( .D(ID_EX__n35), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[7]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_6_ ( .D(ID_EX__n50), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[6]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_5_ ( .D(ID_EX__n1), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[5]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_4_ ( .D(ID_EX__n26), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[4]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_3_ ( .D(ID_EX__n2), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[3]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_2_ ( .D(ID_EX__n217), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[2]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_1_ ( .D(ID_EX__n22), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[1]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___imm_out_reg_0_ ( .D(ID_EX__n179), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_imm[0]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_31_ ( .D(ID_EX__n348), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n810) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_30_ ( .D(ID_EX__n314), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n811) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_29_ ( .D(ID_EX__n460), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n812) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_28_ ( .D(ID_EX__n546), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n813) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_27_ ( .D(ID_EX__n279), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n814) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_26_ ( .D(ID_EX__n461), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n815) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_25_ ( .D(ID_EX__n547), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n816) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_24_ ( .D(ID_EX__n184), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_24_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_23_ ( .D(ID_EX__n349), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_23_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_22_ ( .D(ID_EX__n376), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_22_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_21_ ( .D(ID_EX__n548), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_21_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_20_ ( .D(ID_EX__n341), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_20_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_19_ ( .D(ID_EX__n462), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_19_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_18_ ( .D(ID_EX__n550), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_18_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_17_ ( .D(ID_EX__n350), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_17_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_16_ ( .D(ID_EX__n377), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_16_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_15_ ( .D(ID_EX__n551), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_15_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_14_ ( .D(ID_EX__n256), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n817) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_13_ ( .D(ID_EX__n227), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n818) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_12_ ( .D(ID_EX__n549), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n819) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_11_ ( .D(ID_EX__n351), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_11_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_10_ ( .D(ID_EX__n378), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_10_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_9_ ( .D(ID_EX__n431), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_9_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_8_ ( .D(ID_EX__n379), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_8_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_7_ ( .D(ID_EX__n432), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_inst_7_) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_6_ ( .D(ID_EX__n385), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n820) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_5_ ( .D(ID_EX__n232), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n821) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_4_ ( .D(ID_EX__n433), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n822) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_3_ ( .D(ID_EX__n410), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n823) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_2_ ( .D(ID_EX__n552), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n824) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_1_ ( .D(ID_EX__n369), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n825) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_out_reg_0_ ( .D(ID_EX__n406), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n826) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_31_ ( .D(ID_EX__n315), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX__n827) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_30_ ( .D(ID_EX__n342), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX__n828) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_29_ ( .D(ID_EX__n352), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX__n829) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_28_ ( .D(ID_EX__n257), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[28]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_27_ ( .D(ID_EX__n320), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[27]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_26_ ( .D(ID_EX__n316), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[26]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_25_ ( .D(ID_EX__n380), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[25]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_24_ ( .D(ID_EX__n343), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX__n830) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_23_ ( .D(ID_EX__n321), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX__n831) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_22_ ( .D(ID_EX__n353), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[22]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_21_ ( .D(ID_EX__n281), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[21]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_20_ ( .D(ID_EX__n228), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[20]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_19_ ( .D(ID_EX__n344), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX__n832) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_18_ ( .D(ID_EX__n381), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[18]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_17_ ( .D(ID_EX__n282), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[17]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_16_ ( .D(ID_EX__n259), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[16]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_15_ ( .D(ID_EX__n382), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[15]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_14_ ( .D(ID_EX__n230), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[14]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_13_ ( .D(ID_EX__n383), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[13]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_12_ ( .D(ID_EX__n322), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[12]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_11_ ( .D(ID_EX__n434), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX__n833) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_10_ ( .D(ID_EX__n323), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[10]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_9_ ( .D(ID_EX__n231), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[9]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_8_ ( .D(ID_EX__n283), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[8]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_7_ ( .D(ID_EX__n324), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[7]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_6_ ( .D(ID_EX__n225), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[6]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_5_ ( .D(ID_EX__n384), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[5]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_4_ ( .D(ID_EX__n284), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX__n834) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_3_ ( .D(ID_EX__n229), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[3]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_2_ ( .D(ID_EX__n345), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[2]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_1_ ( .D(ID_EX__n280), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[1]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___inst_addr_out_reg_0_ ( .D(ID_EX__n317), .CLK(clk), .SETN(
        n361), .RESETN(ID_EX__n569), .QN(ID_EX_inst_addr[0]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rd_out_reg_4_ ( .D(ID_EX__n318), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n835) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rd_out_reg_3_ ( .D(ID_EX__n346), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_rd[3]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rd_out_reg_2_ ( .D(ID_EX__n375), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_rd[2]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rd_out_reg_1_ ( .D(ID_EX__n319), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n836) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rd_out_reg_0_ ( .D(ID_EX__n347), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_rd[0]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rs1_out_reg_4_ ( .D(ID_EX__n307), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_rs1[4]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rs1_out_reg_3_ ( .D(ID_EX__n467), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_rs1[3]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rs1_out_reg_2_ ( .D(ID_EX__n370), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n837) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rs1_out_reg_1_ ( .D(ID_EX__n337), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n838) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rs1_out_reg_0_ ( .D(ID_EX__n278), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n839) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rs2_out_reg_4_ ( .D(ID_EX__n153), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_rs2[4]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rs2_out_reg_3_ ( .D(ID_EX__n325), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_rs2[3]) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rs2_out_reg_2_ ( .D(ID_EX__n183), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n840) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rs2_out_reg_1_ ( .D(ID_EX__n557), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n841) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___rs2_out_reg_0_ ( .D(ID_EX__n466), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n842) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___Branch_out_reg ( .D(ID_EX__n3), .CLK(clk), .SETN(ID_EX__ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX_Branch) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___MemRead_out_reg ( .D(ID_EX__n53), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n735) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___MemtoReg_out_reg ( .D(ID_EX__n313), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n736) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___MemWrite_out_reg ( .D(ID_EX__n226), .CLK(clk), .SETN(ID_EX__n361), 
        .RESETN(ID_EX__n569), .QN(ID_EX__n737) );
  CKINVDCx10_ASAP7_75t_R ID_EX___U363 ( .A(rst), .Y(ID_EX__n361) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_0_ ( .D(ID_EX__n9), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n771) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_16_ ( .D(ID_EX__n19), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n755) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_6_ ( .D(ID_EX__n15), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n765) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_25_ ( .D(ID_EX__n69), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n746) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_8_ ( .D(ID_EX__n61), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n763) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_3_ ( .D(ID_EX__n51), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n768) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_21_ ( .D(ID_EX__n56), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__ID_EX__n569), .QN(ID_EX__n750) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_20_ ( .D(ID_EX__n66), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n751) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_18_ ( .D(ID_EX__n59), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n753) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_4_ ( .D(ID_EX__n65), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n767) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_2_ ( .D(ID_EX__n25), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n769) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_22_ ( .D(ID_EX__n75), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n749) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_1_ ( .D(ID_EX__n47), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n770) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_5_ ( .D(ID_EX__n4), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n766) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_11_ ( .D(ID_EX__n12), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n760) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_11_ ( .D(ID_EX__n8), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n792) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_13_ ( .D(ID_EX__n54), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n758) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_13_ ( .D(ID_EX__n72), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n790) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_10_ ( .D(ID_EX__n18), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n761) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_17_ ( .D(ID_EX__n55), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n754) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_10_ ( .D(ID_EX__n10), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n793) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_9_ ( .D(ID_EX__n28), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n762) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_7_ ( .D(ID_EX__n39), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n796) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_30_ ( .D(ID_EX__n63), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n741) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_31_ ( .D(ID_EX__n36), .CLK(clk), 
        .SETN(ID_EX__ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n740) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_7_ ( .D(ID_EX__n31), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n764) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_9_ ( .D(ID_EX__n30), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n794) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_24_ ( .D(ID_EX__n11), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n747) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_15_ ( .D(ID_EX__n52), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n756) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_19_ ( .D(ID_EX__n58), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n752) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_23_ ( .D(ID_EX__n73), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n748) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_12_ ( .D(ID_EX__n74), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n759) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_17_ ( .D(ID_EX__n37), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n786) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_14_ ( .D(ID_EX__n29), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n789) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_31_ ( .D(ID_EX__n40), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n772) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_28_ ( .D(ID_EX__n42), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n775) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_14_ ( .D(ID_EX__n16), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n757) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_24_ ( .D(ID_EX__n49), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n779) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_15_ ( .D(ID_EX__n7), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__ID_EX__n788) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_19_ ( .D(ID_EX__n23), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n784) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_28_ ( .D(ID_EX__n62), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n743) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_26_ ( .D(ID_EX__n34), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n777) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_26_ ( .D(ID_EX__n20), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n745) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_27_ ( .D(ID_EX__n21), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n776) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_30_ ( .D(ID_EX__n70), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n773) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_29_ ( .D(ID_EX__n6), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n774) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_27_ ( .D(ID_EX__n57), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n744) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_1_out_reg_29_ ( .D(ID_EX__n60), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n742) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_23_ ( .D(ID_EX__n44), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n780) );
  DFFASRHQNx1_ASAP7_75t_R ID_EX___read_reg_data_2_out_reg_12_ ( .D(ID_EX__n27), .CLK(clk), 
        .SETN(ID_EX__n361), .RESETN(ID_EX__n569), .QN(ID_EX__n791) );
  TIEHIx1_ASAP7_75t_R ID_EX___U3 ( .H(ID_EX__n569) );
  NAND2xp5_ASAP7_75t_R ID_EX___U4 ( .A(ID_EX__n594), .B(ID_read_reg_data_1[9]), .Y(ID_EX__n28) );
  NAND2xp5_ASAP7_75t_R ID_EX___U5 ( .A(ID_EX__n592), .B(ID_read_reg_data_2[21]), .Y(ID_EX__n33) );
  NAND2xp67_ASAP7_75t_R ID_EX___U6 ( .A(ID_EX__n581), .B(ID_read_reg_data_2[15]), .Y(ID_EX__n7) );
  BUFx2_ASAP7_75t_R ID_EX___U7 ( .A(ID_EX__n831), .Y(ID_EX__n481) );
  BUFx6f_ASAP7_75t_R ID_EX___U8 ( .A(ID_EX__n481), .Y(ID_EX_inst_addr[23]) );
  NAND2xp5_ASAP7_75t_R ID_EX___U9 ( .A(ID_EX__n599), .B(ID_read_reg_data_1[6]), .Y(ID_EX__n15) );
  NAND2xp5_ASAP7_75t_R ID_EX___U10 ( .A(ID_EX__n582), .B(ID_read_reg_data_2[25]), .Y(ID_EX__n14) );
  INVx1_ASAP7_75t_R ID_EX___U11 ( .A(ID_EX__n713), .Y(ID_EX__n1) );
  NAND2xp5_ASAP7_75t_R ID_EX___U12 ( .A(ID_EX__n158), .B(ID_read_reg_data_2[24]), .Y(ID_EX__n49) );
  NAND2xp5_ASAP7_75t_R ID_EX___U13 ( .A(ID_imm[3]), .B(ID_EX__n584), .Y(ID_EX__n2) );
  INVx1_ASAP7_75t_R ID_EX___U14 ( .A(ID_EX__n641), .Y(ID_EX__n177) );
  BUFx3_ASAP7_75t_R ID_EX___U15 ( .A(ID_EX__n830), .Y(ID_EX_inst_addr[24]) );
  BUFx3_ASAP7_75t_R ID_EX___U16 ( .A(ID_EX__n833), .Y(ID_EX_inst_addr[11]) );
  NAND2xp5_ASAP7_75t_R ID_EX___U17 ( .A(ID_EX__n583), .B(ID_read_reg_data_2[26]), .Y(ID_EX__n34) );
  INVx1_ASAP7_75t_R ID_EX___U18 ( .A(ID_EX__n681), .Y(ID_EX__n217) );
  NAND2xp5_ASAP7_75t_R ID_EX___U19 ( .A(ID_EX__n575), .B(ID_Branch), .Y(ID_EX__n3) );
  BUFx3_ASAP7_75t_R ID_EX___U20 ( .A(ID_EX__n640), .Y(ID_EX__n182) );
  NAND2xp5_ASAP7_75t_R ID_EX___U21 ( .A(ID_EX__n116), .B(ID_read_reg_data_1[5]), .Y(ID_EX__n4) );
  NAND2xp5_ASAP7_75t_R ID_EX___U22 ( .A(ID_EX__n115), .B(ID_RegWrite), .Y(ID_EX__n5) );
  INVxp67_ASAP7_75t_R ID_EX___U23 ( .A(ID_EX__n156), .Y(ID_EX__n218) );
  HB1xp67_ASAP7_75t_R ID_EX___U24 ( .A(ID_EX__n644), .Y(ID_EX__n156) );
  NAND2xp5_ASAP7_75t_R ID_EX___U25 ( .A(ID_EX__n606), .B(ID_read_reg_data_1[23]), .Y(ID_EX__n73) );
  NAND2xp5_ASAP7_75t_R ID_EX___U26 ( .A(ID_EX__n581), .B(ID_read_reg_data_2[29]), .Y(ID_EX__n6) );
  NAND2xp5_ASAP7_75t_R ID_EX___U27 ( .A(ID_EX__n590), .B(ID_read_reg_data_2[11]), .Y(ID_EX__n8) );
  NAND2xp5_ASAP7_75t_R ID_EX___U28 ( .A(ID_EX__n593), .B(ID_read_reg_data_1[0]), .Y(ID_EX__n9) );
  NAND2xp5_ASAP7_75t_R ID_EX___U29 ( .A(ID_EX__n590), .B(ID_read_reg_data_2[10]), .Y(ID_EX__n10) );
  BUFx3_ASAP7_75t_R ID_EX___U30 ( .A(ID_EX__n834), .Y(ID_EX_inst_addr[4]) );
  NAND2xp5_ASAP7_75t_R ID_EX___U31 ( .A(ID_EX__n603), .B(ID_read_reg_data_1[24]), .Y(ID_EX__n11) );
  NAND2xp5_ASAP7_75t_R ID_EX___U32 ( .A(ID_EX__n114), .B(ID_read_reg_data_1[11]), .Y(ID_EX__n12) );
  INVx1_ASAP7_75t_R ID_EX___U33 ( .A(ID_EX__n643), .Y(ID_EX__n13) );
  NAND2xp5_ASAP7_75t_R ID_EX___U34 ( .A(ID_EX__n609), .B(ID_read_reg_data_2[2]), .Y(ID_EX__n71) );
  NAND2xp5_ASAP7_75t_R ID_EX___U35 ( .A(ID_EX__n595), .B(ID_read_reg_data_1[14]), .Y(ID_EX__n16) );
  BUFx6f_ASAP7_75t_R ID_EX___U36 ( .A(ID_EX__n477), .Y(ID_EX_rd[4]) );
  INVx1_ASAP7_75t_R ID_EX___U37 ( .A(ID_EX__n663), .Y(ID_EX__n17) );
  BUFx6f_ASAP7_75t_R ID_EX___U38 ( .A(ID_EX__n479), .Y(ID_EX_rd[1]) );
  NAND2xp5_ASAP7_75t_R ID_EX___U39 ( .A(ID_EX__n618), .B(ID_read_reg_data_1[12]), .Y(ID_EX__n74) );
  NAND2xp5_ASAP7_75t_R ID_EX___U40 ( .A(ID_EX__n620), .B(ID_read_reg_data_1[10]), .Y(ID_EX__n18) );
  NAND2xp5_ASAP7_75t_R ID_EX___U41 ( .A(ID_EX__n587), .B(ID_imm[18]), .Y(ID_EX__n24) );
  NAND2xp5_ASAP7_75t_R ID_EX___U42 ( .A(ID_EX__n596), .B(ID_read_reg_data_1[16]), .Y(ID_EX__n19) );
  NAND2xp5_ASAP7_75t_R ID_EX___U43 ( .A(ID_EX__n607), .B(ID_read_reg_data_1[26]), .Y(ID_EX__n20) );
  BUFx3_ASAP7_75t_R ID_EX___U44 ( .A(ID_EX__n808), .Y(ID_EX_imm[15]) );
  NAND2xp5_ASAP7_75t_R ID_EX___U45 ( .A(ID_EX__n157), .B(ID_read_reg_data_2[27]), .Y(ID_EX__n21) );
  INVx1_ASAP7_75t_R ID_EX___U46 ( .A(ID_EX__n670), .Y(ID_EX__n22) );
  NAND2xp5_ASAP7_75t_R ID_EX___U47 ( .A(ID_EX__n576), .B(ID_read_reg_data_2[16]), .Y(ID_EX__n41) );
  NAND2xp5_ASAP7_75t_R ID_EX___U48 ( .A(ID_EX__n619), .B(ID_read_reg_data_2[19]), .Y(ID_EX__n23) );
  NAND2xp5_ASAP7_75t_R ID_EX___U49 ( .A(ID_EX__n580), .B(ID_read_reg_data_1[2]), .Y(ID_EX__n25) );
  INVx1_ASAP7_75t_R ID_EX___U50 ( .A(ID_EX__n702), .Y(ID_EX__n26) );
  NAND2xp5_ASAP7_75t_R ID_EX___U51 ( .A(ID_EX__n591), .B(ID_read_reg_data_2[12]), .Y(ID_EX__n27) );
  INVx2_ASAP7_75t_R ID_EX___U52 ( .A(ID_EX__n148), .Y(ID_EX__n258) );
  BUFx3_ASAP7_75t_R ID_EX___U53 ( .A(ID_EX__n634), .Y(ID_EX__n148) );
  NAND2xp5_ASAP7_75t_R ID_EX___U54 ( .A(ID_EX__n591), .B(ID_read_reg_data_2[14]), .Y(ID_EX__n29) );
  NAND2xp5_ASAP7_75t_R ID_EX___U55 ( .A(ID_EX__n590), .B(ID_read_reg_data_2[9]), .Y(ID_EX__n30) );
  NAND2xp5_ASAP7_75t_R ID_EX___U56 ( .A(ID_EX__n594), .B(ID_read_reg_data_1[7]), .Y(ID_EX__n31) );
  NAND2xp5_ASAP7_75t_R ID_EX___U57 ( .A(ID_EX__n589), .B(ID_read_reg_data_2[4]), .Y(ID_EX__n32) );
  NAND2xp5_ASAP7_75t_R ID_EX___U58 ( .A(ID_EX__n597), .B(ID_read_reg_data_1[21]), .Y(ID_EX__n56) );
  NAND2x1_ASAP7_75t_R ID_EX___U59 ( .A(ID_imm[7]), .B(ID_EX__n585), .Y(ID_EX__n35) );
  NAND2xp5_ASAP7_75t_R ID_EX___U60 ( .A(ID_EX__n621), .B(ID_read_reg_data_1[31]), .Y(ID_EX__n36) );
  NAND2xp5_ASAP7_75t_R ID_EX___U61 ( .A(ID_EX__n610), .B(ID_read_reg_data_2[17]), .Y(ID_EX__n37) );
  NAND2xp5_ASAP7_75t_R ID_EX___U62 ( .A(ID_EX__n602), .B(ID_read_reg_data_2[1]), .Y(ID_EX__n38) );
  BUFx3_ASAP7_75t_R ID_EX___U63 ( .A(ID_EX__n809), .Y(ID_EX_imm[11]) );
  NAND2xp5_ASAP7_75t_R ID_EX___U64 ( .A(ID_EX__n594), .B(ID_read_reg_data_2[7]), .Y(ID_EX__n39) );
  NAND2xp5_ASAP7_75t_R ID_EX___U65 ( .A(ID_EX__n593), .B(ID_read_reg_data_2[31]), .Y(ID_EX__n40) );
  NAND2xp5_ASAP7_75t_R ID_EX___U66 ( .A(ID_EX__n587), .B(ID_read_reg_data_2[28]), .Y(ID_EX__n42) );
  NAND2xp5_ASAP7_75t_R ID_EX___U67 ( .A(ID_EX__n572), .B(ID_read_reg_data_2[18]), .Y(ID_EX__n43) );
  NAND2xp5_ASAP7_75t_R ID_EX___U68 ( .A(ID_EX__n592), .B(ID_read_reg_data_2[23]), .Y(ID_EX__n44) );
  NAND2xp5_ASAP7_75t_R ID_EX___U69 ( .A(ID_EX__n575), .B(ID_read_reg_data_2[20]), .Y(ID_EX__n45) );
  NAND2xp5_ASAP7_75t_R ID_EX___U70 ( .A(ID_EX__n592), .B(ID_read_reg_data_2[22]), .Y(ID_EX__n46) );
  NAND2xp5_ASAP7_75t_R ID_EX___U71 ( .A(ID_EX__n615), .B(ID_read_reg_data_1[1]), .Y(ID_EX__n47) );
  NAND2xp5_ASAP7_75t_R ID_EX___U72 ( .A(ID_EX__n591), .B(ID_read_reg_data_2[13]), .Y(ID_EX__n72) );
  NAND2xp5_ASAP7_75t_R ID_EX___U73 ( .A(ID_EX__n589), .B(ID_read_reg_data_2[3]), .Y(ID_EX__n48) );
  NAND2xp5_ASAP7_75t_R ID_EX___U74 ( .A(ID_EX__n597), .B(ID_read_reg_data_1[20]), .Y(ID_EX__n66) );
  INVx1_ASAP7_75t_R ID_EX___U75 ( .A(ID_EX__n724), .Y(ID_EX__n50) );
  NAND2xp5_ASAP7_75t_R ID_EX___U76 ( .A(ID_EX__n596), .B(ID_read_reg_data_1[17]), .Y(ID_EX__n55) );
  NAND2xp5_ASAP7_75t_R ID_EX___U77 ( .A(ID_EX__n594), .B(ID_read_reg_data_1[3]), .Y(ID_EX__n51) );
  NAND2xp5_ASAP7_75t_R ID_EX___U78 ( .A(ID_EX__n614), .B(ID_read_reg_data_1[22]), .Y(ID_EX__n75) );
  INVx1_ASAP7_75t_R ID_EX___U79 ( .A(ID_EX__n639), .Y(ID_EX__n313) );
  NAND2xp5_ASAP7_75t_R ID_EX___U80 ( .A(ID_EX__n595), .B(ID_read_reg_data_1[15]), .Y(ID_EX__n52) );
  BUFx3_ASAP7_75t_R ID_EX___U81 ( .A(ID_EX__n835), .Y(ID_EX__n477) );
  NAND2xp5_ASAP7_75t_R ID_EX___U82 ( .A(ID_EX__n121), .B(ID_MemRead), .Y(ID_EX__n53) );
  NAND2xp5_ASAP7_75t_R ID_EX___U83 ( .A(ID_EX__n597), .B(ID_read_reg_data_1[19]), .Y(ID_EX__n58) );
  BUFx3_ASAP7_75t_R ID_EX___U84 ( .A(ID_EX__n836), .Y(ID_EX__n479) );
  NAND2xp5_ASAP7_75t_R ID_EX___U85 ( .A(ID_EX__n595), .B(ID_read_reg_data_1[13]), .Y(ID_EX__n54) );
  NAND2xp5_ASAP7_75t_R ID_EX___U86 ( .A(ID_EX__n157), .B(ID_read_reg_data_1[27]), .Y(ID_EX__n57) );
  NAND2xp5_ASAP7_75t_R ID_EX___U87 ( .A(ID_EX__ID_EX__n596), .B(ID_read_reg_data_1[18]), .Y(ID_EX__n59) );
  NAND2xp5_ASAP7_75t_R ID_EX___U88 ( .A(ID_EX__n598), .B(ID_read_reg_data_1[29]), .Y(ID_EX__n60) );
  NAND2xp5_ASAP7_75t_R ID_EX___U89 ( .A(ID_EX__n594), .B(ID_read_reg_data_1[8]), .Y(ID_EX__n61) );
  NAND2xp5_ASAP7_75t_R ID_EX___U90 ( .A(ID_EX__n618), .B(ID_read_reg_data_1[28]), .Y(ID_EX__n62) );
  NAND2xp5_ASAP7_75t_R ID_EX___U91 ( .A(ID_EX__n598), .B(ID_read_reg_data_1[30]), .Y(ID_EX__n63) );
  NAND2xp5_ASAP7_75t_R ID_EX___U92 ( .A(ID_EX__n605), .B(ID_read_reg_data_2[8]), .Y(ID_EX__n64) );
  NAND2xp5_ASAP7_75t_R ID_EX___U93 ( .A(ID_EX__n602), .B(ID_read_reg_data_1[4]), .Y(ID_EX__n65) );
  NAND2xp5_ASAP7_75t_R ID_EX___U94 ( .A(ID_EX__n609), .B(ID_read_reg_data_2[0]), .Y(ID_EX__n67) );
  AND2x2_ASAP7_75t_R ID_EX___U95 ( .A(n40), .B(ID_EX__n570), .Y(ID_EX__n636) );
  NAND2xp5_ASAP7_75t_R ID_EX___U96 ( .A(ID_EX__n580), .B(ID_read_reg_data_2[6]), .Y(ID_EX__n68) );
  NAND2xp5_ASAP7_75t_R ID_EX___U97 ( .A(ID_EX__n610), .B(ID_read_reg_data_1[25]), .Y(ID_EX__n69) );
  NAND2xp5_ASAP7_75t_R ID_EX___U98 ( .A(ID_EX__n593), .B(ID_read_reg_data_2[30]), .Y(ID_EX__n70) );
  NAND2xp5_ASAP7_75t_R ID_EX___U99 ( .A(ID_EX__n589), .B(ID_read_reg_data_2[5]), .Y(ID_EX__n76) );
  AND2x2_ASAP7_75t_R ID_EX___U100 ( .A(n30), .B(ID_EX__n572), .Y(ID_EX__n629) );
  AND2x2_ASAP7_75t_R ID_EX___U101 ( .A(n43), .B(ID_EX__n570), .Y(ID_EX__n633) );
  BUFx3_ASAP7_75t_R ID_EX___U102 ( .A(ID_EX__n653), .Y(ID_EX__n88) );
  BUFx3_ASAP7_75t_R ID_EX___U103 ( .A(ID_EX__n652), .Y(ID_EX__n90) );
  AND2x2_ASAP7_75t_R ID_EX___U104 ( .A(n26), .B(ID_EX__n571), .Y(ID_EX__n638) );
  AND2x2_ASAP7_75t_R ID_EX___U105 ( .A(n45), .B(ID_EX__n571), .Y(ID_EX__n628) );
  BUFx2_ASAP7_75t_R ID_EX___U106 ( .A(ID_EX__n664), .Y(ID_EX__n77) );
  BUFx2_ASAP7_75t_R ID_EX___U107 ( .A(ID_EX__n662), .Y(ID_EX__n78) );
  BUFx2_ASAP7_75t_R ID_EX___U108 ( .A(ID_EX__n661), .Y(ID_EX__n79) );
  BUFx2_ASAP7_75t_R ID_EX___U109 ( .A(ID_EX__n660), .Y(ID_EX__n80) );
  BUFx2_ASAP7_75t_R ID_EX___U110 ( .A(ID_EX__n658), .Y(ID_EX__n81) );
  BUFx2_ASAP7_75t_R ID_EX___U111 ( .A(ID_EX__n657), .Y(ID_EX__n82) );
  BUFx2_ASAP7_75t_R ID_EX___U112 ( .A(ID_EX__n656), .Y(ID_EX__n83) );
  BUFx2_ASAP7_75t_R ID_EX___U113 ( .A(ID_EX__n655), .Y(ID_EX__n84) );
  BUFx2_ASAP7_75t_R ID_EX___U114 ( .A(ID_EX__n651), .Y(ID_EX__n85) );
  BUFx2_ASAP7_75t_R ID_EX___U115 ( .A(ID_EX__n654), .Y(ID_EX__n86) );
  BUFx2_ASAP7_75t_R ID_EX___U116 ( .A(ID_EX__n650), .Y(ID_EX__n87) );
  BUFx2_ASAP7_75t_R ID_EX___U117 ( .A(ID_EX__n649), .Y(ID_EX__n89) );
  BUFx2_ASAP7_75t_R ID_EX___U118 ( .A(ID_EX__n648), .Y(ID_EX__n91) );
  BUFx12f_ASAP7_75t_R ID_EX___U119 ( .A(ID_EX__n120), .Y(ID_EX__n92) );
  BUFx12f_ASAP7_75t_R ID_EX___U120 ( .A(ID_EX__n92), .Y(ID_EX__n93) );
  BUFx12f_ASAP7_75t_R ID_EX___U121 ( .A(ID_EX__n122), .Y(ID_EX__n94) );
  BUFx12f_ASAP7_75t_R ID_EX___U122 ( .A(ID_EX__n105), .Y(ID_EX__n95) );
  BUFx12f_ASAP7_75t_R ID_EX___U123 ( .A(ID_EX__n105), .Y(ID_EX__n96) );
  BUFx12f_ASAP7_75t_R ID_EX___U124 ( .A(ID_EX__n106), .Y(ID_EX__n97) );
  BUFx12f_ASAP7_75t_R ID_EX___U125 ( .A(ID_EX__n107), .Y(ID_EX__n98) );
  BUFx12f_ASAP7_75t_R ID_EX___U126 ( .A(ID_EX__n98), .Y(ID_EX__n99) );
  BUFx12f_ASAP7_75t_R ID_EX___U127 ( .A(ID_EX__n108), .Y(ID_EX__n100) );
  BUFx12f_ASAP7_75t_R ID_EX___U128 ( .A(ID_EX__n109), .Y(ID_EX__n101) );
  BUFx12f_ASAP7_75t_R ID_EX___U129 ( .A(ID_EX__n101), .Y(ID_EX__n102) );
  BUFx12f_ASAP7_75t_R ID_EX___U130 ( .A(ID_EX__n104), .Y(ID_EX__n103) );
  BUFx12f_ASAP7_75t_R ID_EX___U131 ( .A(ID_EX__n110), .Y(ID_EX__n104) );
  BUFx12f_ASAP7_75t_R ID_EX___U132 ( .A(ID_EX__n112), .Y(ID_EX__n105) );
  BUFx12f_ASAP7_75t_R ID_EX___U133 ( .A(ID_EX__n113), .Y(ID_EX__n106) );
  BUFx12f_ASAP7_75t_R ID_EX___U134 ( .A(ID_EX__n111), .Y(ID_EX__n107) );
  BUFx12f_ASAP7_75t_R ID_EX___U135 ( .A(ID_EX__n119), .Y(ID_EX__n108) );
  BUFx12f_ASAP7_75t_R ID_EX___U136 ( .A(ID_EX__n118), .Y(ID_EX__n109) );
  BUFx12f_ASAP7_75t_R ID_EX___U137 ( .A(ID_EX__n117), .Y(ID_EX__n110) );
  BUFx12f_ASAP7_75t_R ID_EX___U138 ( .A(ID_EX__n115), .Y(ID_EX__n111) );
  BUFx12f_ASAP7_75t_R ID_EX___U139 ( .A(ID_EX__n116), .Y(ID_EX__n112) );
  BUFx12f_ASAP7_75t_R ID_EX___U140 ( .A(ID_EX__n121), .Y(ID_EX__n113) );
  BUFx12f_ASAP7_75t_R ID_EX___U141 ( .A(ID_EX__n99), .Y(ID_EX__n114) );
  BUFx12f_ASAP7_75t_R ID_EX___U142 ( .A(ID_EX__n620), .Y(ID_EX__n115) );
  BUFx12f_ASAP7_75t_R ID_EX___U143 ( .A(ID_EX__n618), .Y(ID_EX__n116) );
  BUFx12f_ASAP7_75t_R ID_EX___U144 ( .A(ID_EX__n617), .Y(ID_EX__n117) );
  BUFx12f_ASAP7_75t_R ID_EX___U145 ( .A(ID_EX__n616), .Y(ID_EX__n118) );
  BUFx12f_ASAP7_75t_R ID_EX___U146 ( .A(ID_EX__n619), .Y(ID_EX__n119) );
  BUFx12f_ASAP7_75t_R ID_EX___U147 ( .A(ID_EX__n622), .Y(ID_EX__n120) );
  BUFx12f_ASAP7_75t_R ID_EX___U148 ( .A(ID_EX__n124), .Y(ID_EX__n121) );
  BUFx12f_ASAP7_75t_R ID_EX___U149 ( .A(ID_EX__n123), .Y(ID_EX__n122) );
  BUFx12f_ASAP7_75t_R ID_EX___U150 ( .A(ID_EX__n127), .Y(ID_EX__n123) );
  BUFx12f_ASAP7_75t_R ID_EX___U151 ( .A(ID_EX__n128), .Y(ID_EX__n124) );
  BUFx12f_ASAP7_75t_R ID_EX___U152 ( .A(ID_EX__n94), .Y(ID_EX__n125) );
  BUFx12f_ASAP7_75t_R ID_EX___U153 ( .A(ID_EX__n94), .Y(ID_EX__n126) );
  BUFx12f_ASAP7_75t_R ID_EX___U154 ( .A(ID_EX__n608), .Y(ID_EX__n127) );
  BUFx12f_ASAP7_75t_R ID_EX___U155 ( .A(ID_EX__n129), .Y(ID_EX__n128) );
  BUFx12f_ASAP7_75t_R ID_EX___U156 ( .A(ID_EX__n604), .Y(ID_EX__n129) );
  BUFx12f_ASAP7_75t_R ID_EX___U157 ( .A(ID_EX__n613), .Y(ID_EX__n570) );
  BUFx2_ASAP7_75t_R ID_EX___U158 ( .A(ID_EX__n647), .Y(ID_EX__n130) );
  AND2x2_ASAP7_75t_R ID_EX___U159 ( .A(ID_imm[31]), .B(ID_EX__n582), .Y(ID_EX__n664) );
  INVx1_ASAP7_75t_R ID_EX___U160 ( .A(ID_EX__n77), .Y(ID_EX__n131) );
  BUFx2_ASAP7_75t_R ID_EX___U161 ( .A(ID_EX__n646), .Y(ID_EX__n132) );
  AND2x2_ASAP7_75t_R ID_EX___U162 ( .A(ID_imm[24]), .B(ID_EX__n576), .Y(ID_EX__n656) );
  INVx1_ASAP7_75t_R ID_EX___U163 ( .A(ID_EX__n83), .Y(ID_EX__n133) );
  AND2x2_ASAP7_75t_R ID_EX___U164 ( .A(ID_imm[23]), .B(ID_EX__n576), .Y(ID_EX__n655) );
  INVx1_ASAP7_75t_R ID_EX___U165 ( .A(ID_EX__n84), .Y(ID_EX__n134) );
  AND2x2_ASAP7_75t_R ID_EX___U166 ( .A(ID_imm[22]), .B(ID_EX__n580), .Y(ID_EX__n654) );
  INVx1_ASAP7_75t_R ID_EX___U167 ( .A(ID_EX__n86), .Y(ID_EX__n135) );
  BUFx2_ASAP7_75t_R ID_EX___U168 ( .A(ID_EX__n645), .Y(ID_EX__n136) );
  AND2x2_ASAP7_75t_R ID_EX___U169 ( .A(ID_imm[21]), .B(ID_EX__n571), .Y(ID_EX__n653) );
  INVx1_ASAP7_75t_R ID_EX___U170 ( .A(ID_EX__n88), .Y(ID_EX__n137) );
  BUFx12f_ASAP7_75t_R ID_EX___U171 ( .A(ID_EX__n615), .Y(ID_EX__n612) );
  BUFx12f_ASAP7_75t_R ID_EX___U172 ( .A(ID_EX__n100), .Y(ID_EX__n601) );
  BUFx12f_ASAP7_75t_R ID_EX___U173 ( .A(ID_EX__n101), .Y(ID_EX__n611) );
  BUFx12f_ASAP7_75t_R ID_EX___U174 ( .A(ID_EX__n140), .Y(ID_EX__n138) );
  BUFx12f_ASAP7_75t_R ID_EX___U175 ( .A(ID_EX__n141), .Y(ID_EX__n139) );
  BUFx12f_ASAP7_75t_R ID_EX___U176 ( .A(ID_EX__n97), .Y(ID_EX__n140) );
  BUFx12f_ASAP7_75t_R ID_EX___U177 ( .A(ID_EX__n97), .Y(ID_EX__n141) );
  BUFx12f_ASAP7_75t_R ID_EX___U178 ( .A(ID_EX__n114), .Y(ID_EX__n604) );
  BUFx12f_ASAP7_75t_R ID_EX___U179 ( .A(ID_EX__n92), .Y(ID_EX__n605) );
  BUFx12f_ASAP7_75t_R ID_EX___U180 ( .A(ID_EX__n95), .Y(ID_EX__n603) );
  AND2x2_ASAP7_75t_R ID_EX___U181 ( .A(ID_imm[20]), .B(ID_EX__n603), .Y(ID_EX__n652) );
  INVx1_ASAP7_75t_R ID_EX___U182 ( .A(ID_EX__n90), .Y(ID_EX__n142) );
  AND2x2_ASAP7_75t_R ID_EX___U183 ( .A(ID_imm[19]), .B(ID_EX__n587), .Y(ID_EX__n651) );
  INVx1_ASAP7_75t_R ID_EX___U184 ( .A(ID_EX__n85), .Y(ID_EX__n143) );
  BUFx2_ASAP7_75t_R ID_EX___U185 ( .A(ID_EX__n642), .Y(ID_EX__n144) );
  AND2x2_ASAP7_75t_R ID_EX___U186 ( .A(ID_imm[29]), .B(ID_EX__n587), .Y(ID_EX__n662) );
  INVx1_ASAP7_75t_R ID_EX___U187 ( .A(ID_EX__n78), .Y(ID_EX__n145) );
  AND2x2_ASAP7_75t_R ID_EX___U188 ( .A(ID_imm[17]), .B(ID_EX__n587), .Y(ID_EX__n650) );
  INVx1_ASAP7_75t_R ID_EX___U189 ( .A(ID_EX__n87), .Y(ID_EX__n146) );
  BUFx2_ASAP7_75t_R ID_EX___U190 ( .A(ID_EX__n715), .Y(ID_EX__n147) );
  BUFx2_ASAP7_75t_R ID_EX___U191 ( .A(ID_EX__n630), .Y(ID_EX__n149) );
  AND2x2_ASAP7_75t_R ID_EX___U192 ( .A(ID_imm[28]), .B(ID_EX__n588), .Y(ID_EX__n661) );
  INVx1_ASAP7_75t_R ID_EX___U193 ( .A(ID_EX__n79), .Y(ID_EX__n150) );
  AND2x2_ASAP7_75t_R ID_EX___U194 ( .A(ID_imm[16]), .B(ID_EX__n107), .Y(ID_EX__n649) );
  INVx1_ASAP7_75t_R ID_EX___U195 ( .A(ID_EX__n89), .Y(ID_EX__n151) );
  BUFx2_ASAP7_75t_R ID_EX___U196 ( .A(ID_EX__n730), .Y(ID_EX__n152) );
  INVx1_ASAP7_75t_R ID_EX___U197 ( .A(ID_EX__n638), .Y(ID_EX__n153) );
  AND2x2_ASAP7_75t_R ID_EX___U198 ( .A(ID_imm[10]), .B(ID_EX__n622), .Y(ID_EX__n643) );
  AND2x2_ASAP7_75t_R ID_EX___U199 ( .A(ID_imm[26]), .B(ID_EX__n588), .Y(ID_EX__n658) );
  INVx1_ASAP7_75t_R ID_EX___U200 ( .A(ID_EX__n81), .Y(ID_EX__n154) );
  AND2x2_ASAP7_75t_R ID_EX___U201 ( .A(ID_imm[14]), .B(ID_EX__n99), .Y(ID_EX__n647) );
  INVx1_ASAP7_75t_R ID_EX___U202 ( .A(ID_EX__n130), .Y(ID_EX__n155) );
  BUFx12f_ASAP7_75t_R ID_EX___U203 ( .A(ID_EX__n93), .Y(ID_EX__n606) );
  BUFx12f_ASAP7_75t_R ID_EX___U204 ( .A(ID_EX__n96), .Y(ID_EX__n607) );
  BUFx12f_ASAP7_75t_R ID_EX___U205 ( .A(ID_EX__n578), .Y(ID_EX__n584) );
  BUFx12f_ASAP7_75t_R ID_EX___U206 ( .A(ID_EX__n595), .Y(ID_EX__n585) );
  BUFx12f_ASAP7_75t_R ID_EX___U207 ( .A(ID_EX__n126), .Y(ID_EX__n157) );
  BUFx12f_ASAP7_75t_R ID_EX___U208 ( .A(ID_EX__n125), .Y(ID_EX__n158) );
  BUFx12f_ASAP7_75t_R ID_EX___U209 ( .A(ID_EX__n98), .Y(ID_EX__n608) );
  BUFx12f_ASAP7_75t_R ID_EX___U210 ( .A(ID_EX__n584), .Y(ID_EX__n586) );
  BUFx12f_ASAP7_75t_R ID_EX___U211 ( .A(ID_EX__n192), .Y(ID_EX__n159) );
  BUFx12f_ASAP7_75t_R ID_EX___U212 ( .A(ID_EX__n103), .Y(ID_EX__n610) );
  BUFx12f_ASAP7_75t_R ID_EX___U213 ( .A(ID_EX__n623), .Y(ID_EX__n618) );
  BUFx2_ASAP7_75t_R ID_EX___U214 ( .A(ID_EX__n814), .Y(ID_EX__n160) );
  BUFx12f_ASAP7_75t_R ID_EX___U215 ( .A(ID_EX__n623), .Y(ID_EX__n620) );
  BUFx16f_ASAP7_75t_R ID_EX___U216 ( .A(ID_EX__n162), .Y(ID_EX__n161) );
  BUFx12f_ASAP7_75t_R ID_EX___U217 ( .A(ID_EX__n159), .Y(ID_EX__n162) );
  BUFx6f_ASAP7_75t_R ID_EX___U218 ( .A(ID_EX__n823), .Y(ID_EX_inst_3_) );
  BUFx2_ASAP7_75t_R ID_EX___U219 ( .A(ID_EX__n815), .Y(ID_EX_inst_26_) );
  BUFx12f_ASAP7_75t_R ID_EX___U220 ( .A(ID_EX__n100), .Y(ID_EX__n602) );
  BUFx12f_ASAP7_75t_R ID_EX___U221 ( .A(ID_EX__n623), .Y(ID_EX__n616) );
  BUFx12f_ASAP7_75t_R ID_EX___U222 ( .A(ID_EX__n102), .Y(ID_EX__n609) );
  BUFx12f_ASAP7_75t_R ID_EX___U223 ( .A(ID_EX__n600), .Y(ID_EX__n615) );
  BUFx12f_ASAP7_75t_R ID_EX___U224 ( .A(ID_EX__n202), .Y(ID_EX_inst_14_) );
  BUFx2_ASAP7_75t_R ID_EX___U225 ( .A(ID_EX__n816), .Y(ID_EX_inst_25_) );
  BUFx12f_ASAP7_75t_R ID_EX___U226 ( .A(ID_EX__n614), .Y(ID_EX__n613) );
  BUFx12f_ASAP7_75t_R ID_EX___U227 ( .A(ID_EX__n621), .Y(ID_EX__n614) );
  BUFx12f_ASAP7_75t_R ID_EX___U228 ( .A(ID_EX__n104), .Y(ID_EX__n621) );
  BUFx2_ASAP7_75t_R ID_EX___U229 ( .A(ID_EX__n810), .Y(ID_EX_inst_31_) );
  BUFx12f_ASAP7_75t_R ID_EX___U230 ( .A(ID_EX__n623), .Y(ID_EX__n619) );
  BUFx12f_ASAP7_75t_R ID_EX___U231 ( .A(ID_EX__n623), .Y(ID_EX__n617) );
  BUFx2_ASAP7_75t_R ID_EX___U232 ( .A(ID_EX__n679), .Y(ID_EX__n168) );
  BUFx2_ASAP7_75t_R ID_EX___U233 ( .A(ID_EX__n668), .Y(ID_EX__n169) );
  BUFx2_ASAP7_75t_R ID_EX___U234 ( .A(ID_EX__n723), .Y(ID_EX__n170) );
  AND2x2_ASAP7_75t_R ID_EX___U235 ( .A(ID_imm[9]), .B(ID_EX__n122), .Y(ID_EX__n642) );
  INVx1_ASAP7_75t_R ID_EX___U236 ( .A(ID_EX__n144), .Y(ID_EX__n171) );
  AND2x4_ASAP7_75t_R ID_EX___U237 ( .A(ID_imm[0]), .B(ID_EX__n583), .Y(ID_EX__n659) );
  BUFx2_ASAP7_75t_R ID_EX___U238 ( .A(ID_EX__n709), .Y(ID_EX__n172) );
  BUFx2_ASAP7_75t_R ID_EX___U239 ( .A(ID_EX__n719), .Y(ID_EX__n173) );
  AND2x2_ASAP7_75t_R ID_EX___U240 ( .A(ID_imm[25]), .B(ID_EX__n613), .Y(ID_EX__n657) );
  INVx1_ASAP7_75t_R ID_EX___U241 ( .A(ID_EX__n82), .Y(ID_EX__n174) );
  AND2x2_ASAP7_75t_R ID_EX___U242 ( .A(ID_imm[15]), .B(ID_EX__n124), .Y(ID_EX__n648) );
  INVx1_ASAP7_75t_R ID_EX___U243 ( .A(ID_EX__n91), .Y(ID_EX__n175) );
  BUFx6f_ASAP7_75t_R ID_EX___U244 ( .A(ID_EX__n216), .Y(ID_EX_rs2[1]) );
  AND2x2_ASAP7_75t_R ID_EX___U245 ( .A(ID_EX__n621), .B(ID_ALUSrc), .Y(ID_EX__n641) );
  AND2x2_ASAP7_75t_R ID_EX___U246 ( .A(ID_imm[4]), .B(ID_EX__n584), .Y(ID_EX__n702) );
  INVx1_ASAP7_75t_R ID_EX___U247 ( .A(ID_EX__n659), .Y(ID_EX__n179) );
  BUFx2_ASAP7_75t_R ID_EX___U248 ( .A(ID_EX__n725), .Y(ID_EX__n180) );
  BUFx2_ASAP7_75t_R ID_EX___U249 ( .A(ID_EX__n704), .Y(ID_EX__n181) );
  INVx1_ASAP7_75t_R ID_EX___U250 ( .A(ID_EX__n636), .Y(ID_EX__n183) );
  AND2x4_ASAP7_75t_R ID_EX___U251 ( .A(IF_ID_inst[24]), .B(ID_EX__n600), .Y(ID_EX__n691) );
  INVx1_ASAP7_75t_R ID_EX___U252 ( .A(ID_EX__n691), .Y(ID_EX__n184) );
  AND2x2_ASAP7_75t_R ID_EX___U253 ( .A(ID_imm[13]), .B(ID_EX__n586), .Y(ID_EX__n646) );
  INVx1_ASAP7_75t_R ID_EX___U254 ( .A(ID_EX__n132), .Y(ID_EX__n185) );
  BUFx2_ASAP7_75t_R ID_EX___U255 ( .A(ID_EX__n785), .Y(ID_EX__n186) );
  BUFx2_ASAP7_75t_R ID_EX___U256 ( .A(ID_EX__n160), .Y(ID_EX_inst_27_) );
  BUFx3_ASAP7_75t_R ID_EX___U257 ( .A(ID_EX__n189), .Y(ID_EX__n188) );
  BUFx2_ASAP7_75t_R ID_EX___U258 ( .A(ID_EX__n820), .Y(ID_EX__n189) );
  BUFx3_ASAP7_75t_R ID_EX___U259 ( .A(ID_EX__n191), .Y(ID_EX_MemRead) );
  BUFx2_ASAP7_75t_R ID_EX___U260 ( .A(ID_EX__n735), .Y(ID_EX__n191) );
  BUFx12_ASAP7_75t_R ID_EX___U261 ( .A(ID_EX__n738), .Y(ID_EX__n192) );
  CKINVDCx20_ASAP7_75t_R ID_EX___U262 ( .A(ID_EX__n161), .Y(ID_EX__n193) );
  CKINVDCx20_ASAP7_75t_R ID_EX___U263 ( .A(ID_EX__n193), .Y(ID_EX_ALUSrc) );
  BUFx6f_ASAP7_75t_R ID_EX___U264 ( .A(ID_EX__n242), .Y(ID_EX_rs2[0]) );
  BUFx2_ASAP7_75t_R ID_EX___U265 ( .A(ID_EX__n772), .Y(ID_EX__n196) );
  BUFx12f_ASAP7_75t_R ID_EX___U266 ( .A(ID_EX__n562), .Y(ID_EX_inst_13_) );
  BUFx3_ASAP7_75t_R ID_EX___U267 ( .A(ID_EX__n199), .Y(ID_EX__n198) );
  BUFx2_ASAP7_75t_R ID_EX___U268 ( .A(ID_EX__n804), .Y(ID_EX__n199) );
  BUFx3_ASAP7_75t_R ID_EX___U269 ( .A(ID_EX__n201), .Y(ID_EX__n200) );
  BUFx2_ASAP7_75t_R ID_EX___U270 ( .A(ID_EX__n821), .Y(ID_EX__n201) );
  BUFx12f_ASAP7_75t_R ID_EX___U271 ( .A(ID_EX__n623), .Y(ID_EX__n622) );
  CKINVDCx20_ASAP7_75t_R ID_EX___U272 ( .A(ID_flush), .Y(ID_EX__n623) );
  BUFx12f_ASAP7_75t_R ID_EX___U273 ( .A(ID_EX__n203), .Y(ID_EX__n202) );
  BUFx12f_ASAP7_75t_R ID_EX___U274 ( .A(ID_EX__n411), .Y(ID_EX__n203) );
  BUFx2_ASAP7_75t_R ID_EX___U275 ( .A(ID_EX__n678), .Y(ID_EX__n204) );
  BUFx2_ASAP7_75t_R ID_EX___U276 ( .A(ID_EX__n671), .Y(ID_EX__n205) );
  BUFx2_ASAP7_75t_R ID_EX___U277 ( .A(ID_EX__n731), .Y(ID_EX__n206) );
  BUFx2_ASAP7_75t_R ID_EX___U278 ( .A(ID_EX__n708), .Y(ID_EX__n207) );
  BUFx2_ASAP7_75t_R ID_EX___U279 ( .A(ID_EX__n624), .Y(ID_EX__n208) );
  BUFx2_ASAP7_75t_R ID_EX___U280 ( .A(ID_EX__n718), .Y(ID_EX__n209) );
  BUFx2_ASAP7_75t_R ID_EX___U281 ( .A(ID_EX__n712), .Y(ID_EX__n210) );
  AND2x2_ASAP7_75t_R ID_EX___U282 ( .A(ID_imm[27]), .B(ID_EX__n588), .Y(ID_EX__n660) );
  INVx1_ASAP7_75t_R ID_EX___U283 ( .A(ID_EX__n80), .Y(ID_EX__n211) );
  BUFx2_ASAP7_75t_R ID_EX___U284 ( .A(ID_EX__n790), .Y(ID_EX__n212) );
  BUFx2_ASAP7_75t_R ID_EX___U285 ( .A(ID_EX__n779), .Y(ID_EX__n213) );
  BUFx3_ASAP7_75t_R ID_EX___U286 ( .A(ID_EX__n215), .Y(ID_EX__n214) );
  BUFx2_ASAP7_75t_R ID_EX___U287 ( .A(ID_EX__n841), .Y(ID_EX__n215) );
  BUFx6f_ASAP7_75t_R ID_EX___U288 ( .A(ID_EX__n470), .Y(ID_EX__n216) );
  AND2x2_ASAP7_75t_R ID_EX___U289 ( .A(ID_imm[2]), .B(ID_EX__n584), .Y(ID_EX__n681) );
  AND2x2_ASAP7_75t_R ID_EX___U290 ( .A(ID_EX__n586), .B(ID_imm[11]), .Y(ID_EX__n644) );
  BUFx2_ASAP7_75t_R ID_EX___U291 ( .A(ID_EX__n729), .Y(ID_EX__n219) );
  BUFx2_ASAP7_75t_R ID_EX___U292 ( .A(ID_EX__n727), .Y(ID_EX__n220) );
  BUFx2_ASAP7_75t_R ID_EX___U293 ( .A(ID_EX__n722), .Y(ID_EX__n221) );
  BUFx2_ASAP7_75t_R ID_EX___U294 ( .A(ID_EX__n717), .Y(ID_EX__n222) );
  BUFx2_ASAP7_75t_R ID_EX___U295 ( .A(ID_EX__n627), .Y(ID_EX__n223) );
  BUFx2_ASAP7_75t_R ID_EX___U296 ( .A(ID_EX__n632), .Y(ID_EX__n224) );
  AND2x4_ASAP7_75t_R ID_EX___U297 ( .A(IF_ID_inst_addr[6]), .B(ID_EX__n612), .Y(ID_EX__n706) );
  INVx1_ASAP7_75t_R ID_EX___U298 ( .A(ID_EX__n706), .Y(ID_EX__n225) );
  AND2x2_ASAP7_75t_R ID_EX___U299 ( .A(ID_EX__n616), .B(ID_MemWrite), .Y(ID_EX__n640) );
  INVx1_ASAP7_75t_R ID_EX___U300 ( .A(ID_EX__n182), .Y(ID_EX__n226) );
  AND2x2_ASAP7_75t_R ID_EX___U301 ( .A(IF_ID_inst[13]), .B(ID_EX__n140), .Y(ID_EX__n679) );
  INVx1_ASAP7_75t_R ID_EX___U302 ( .A(ID_EX__n168), .Y(ID_EX__n227) );
  AND2x4_ASAP7_75t_R ID_EX___U303 ( .A(IF_ID_inst_addr[20]), .B(ID_EX__n141), .Y(ID_EX__n721) );
  INVx1_ASAP7_75t_R ID_EX___U304 ( .A(ID_EX__n721), .Y(ID_EX__n228) );
  AND2x4_ASAP7_75t_R ID_EX___U305 ( .A(IF_ID_inst_addr[3]), .B(ID_EX__n127), .Y(ID_EX__n703) );
  INVx1_ASAP7_75t_R ID_EX___U306 ( .A(ID_EX__n703), .Y(ID_EX__n229) );
  AND2x2_ASAP7_75t_R ID_EX___U307 ( .A(IF_ID_inst_addr[14]), .B(ID_EX__n575), .Y(ID_EX__n715) );
  INVx1_ASAP7_75t_R ID_EX___U308 ( .A(ID_EX__n147), .Y(ID_EX__n230) );
  AND2x2_ASAP7_75t_R ID_EX___U309 ( .A(IF_ID_inst_addr[9]), .B(ID_EX__n606), .Y(ID_EX__n709) );
  INVx1_ASAP7_75t_R ID_EX___U310 ( .A(ID_EX__n172), .Y(ID_EX__n231) );
  AND2x2_ASAP7_75t_R ID_EX___U311 ( .A(IF_ID_inst[5]), .B(ID_EX__n580), .Y(ID_EX__n671) );
  INVx1_ASAP7_75t_R ID_EX___U312 ( .A(ID_EX__n205), .Y(ID_EX__n232) );
  AND2x2_ASAP7_75t_R ID_EX___U313 ( .A(ID_imm[6]), .B(ID_EX__n585), .Y(ID_EX__n724) );
  BUFx2_ASAP7_75t_R ID_EX___U314 ( .A(ID_EX__n802), .Y(ID_EX__n233) );
  BUFx3_ASAP7_75t_R ID_EX___U315 ( .A(ID_EX__n334), .Y(ID_EX__n234) );
  BUFx4f_ASAP7_75t_R ID_EX___U316 ( .A(ID_EX__n234), .Y(ID_EX__n413) );
  BUFx6f_ASAP7_75t_R ID_EX___U317 ( .A(ID_EX__n300), .Y(ID_EX_inst_addr[31]) );
  BUFx3_ASAP7_75t_R ID_EX___U318 ( .A(ID_EX__n237), .Y(ID_EX__n236) );
  BUFx2_ASAP7_75t_R ID_EX___U319 ( .A(ID_EX__n807), .Y(ID_EX__n237) );
  BUFx3_ASAP7_75t_R ID_EX___U320 ( .A(ID_EX__n239), .Y(ID_EX__n238) );
  BUFx2_ASAP7_75t_R ID_EX___U321 ( .A(ID_EX__n822), .Y(ID_EX__n239) );
  BUFx3_ASAP7_75t_R ID_EX___U322 ( .A(ID_EX__n241), .Y(ID_EX__n240) );
  BUFx2_ASAP7_75t_R ID_EX___U323 ( .A(ID_EX__n842), .Y(ID_EX__n241) );
  BUFx6f_ASAP7_75t_R ID_EX___U324 ( .A(ID_EX__n416), .Y(ID_EX__n242) );
  BUFx12f_ASAP7_75t_R ID_EX___U325 ( .A(ID_EX__n811), .Y(ID_EX__n243) );
  BUFx12f_ASAP7_75t_R ID_EX___U326 ( .A(ID_EX__n374), .Y(ID_EX_imm[19]) );
  BUFx2_ASAP7_75t_R ID_EX___U327 ( .A(ID_EX__n696), .Y(ID_EX__n244) );
  BUFx2_ASAP7_75t_R ID_EX___U328 ( .A(ID_EX__n693), .Y(ID_EX__n245) );
  BUFx2_ASAP7_75t_R ID_EX___U329 ( .A(ID_EX__n686), .Y(ID_EX__n246) );
  BUFx2_ASAP7_75t_R ID_EX___U330 ( .A(ID_EX__n666), .Y(ID_EX__n247) );
  BUFx2_ASAP7_75t_R ID_EX___U331 ( .A(ID_EX__n714), .Y(ID_EX__n248) );
  BUFx2_ASAP7_75t_R ID_EX___U332 ( .A(ID_EX__n711), .Y(ID_EX__n249) );
  BUFx2_ASAP7_75t_R ID_EX___U333 ( .A(ID_EX__n707), .Y(ID_EX__n250) );
  BUFx2_ASAP7_75t_R ID_EX___U334 ( .A(ID_EX__n705), .Y(ID_EX__n251) );
  BUFx2_ASAP7_75t_R ID_EX___U335 ( .A(ID_EX__n626), .Y(ID_EX__n252) );
  BUFx2_ASAP7_75t_R ID_EX___U336 ( .A(ID_EX__n734), .Y(ID_EX__n253) );
  BUFx2_ASAP7_75t_R ID_EX___U337 ( .A(ID_EX__n672), .Y(ID_EX__n254) );
  BUFx2_ASAP7_75t_R ID_EX___U338 ( .A(ID_EX__n637), .Y(ID_EX__n255) );
  AND2x4_ASAP7_75t_R ID_EX___U339 ( .A(IF_ID_inst[14]), .B(ID_EX__n139), .Y(ID_EX__n680) );
  INVx1_ASAP7_75t_R ID_EX___U340 ( .A(ID_EX__n680), .Y(ID_EX__n256) );
  AND2x2_ASAP7_75t_R ID_EX___U341 ( .A(IF_ID_inst_addr[28]), .B(ID_EX__n578), .Y(ID_EX__n730) );
  INVx1_ASAP7_75t_R ID_EX___U342 ( .A(ID_EX__n152), .Y(ID_EX__n257) );
  AND2x2_ASAP7_75t_R ID_EX___U343 ( .A(ID_EX__n123), .B(ID_imm[8]), .Y(ID_EX__n634) );
  AND2x2_ASAP7_75t_R ID_EX___U344 ( .A(ID_imm[5]), .B(ID_EX__n585), .Y(ID_EX__n713) );
  AND2x2_ASAP7_75t_R ID_EX___U345 ( .A(IF_ID_inst_addr[16]), .B(ID_EX__n594), .Y(ID_EX__n717) );
  INVx1_ASAP7_75t_R ID_EX___U346 ( .A(ID_EX__n222), .Y(ID_EX__n259) );
  BUFx2_ASAP7_75t_R ID_EX___U347 ( .A(ID_EX__n261), .Y(ID_EX_RegWrite) );
  BUFx2_ASAP7_75t_R ID_EX___U348 ( .A(ID_EX__n739), .Y(ID_EX__n261) );
  BUFx6f_ASAP7_75t_R ID_EX___U349 ( .A(ID_EX__n303), .Y(ID_EX_rs1[2]) );
  BUFx6f_ASAP7_75t_R ID_EX___U350 ( .A(ID_EX__n306), .Y(ID_EX_rs2[2]) );
  BUFx2_ASAP7_75t_R ID_EX___U351 ( .A(ID_EX__n761), .Y(ID_EX__n264) );
  BUFx2_ASAP7_75t_R ID_EX___U352 ( .A(ID_EX__n794), .Y(ID_EX__n265) );
  BUFx2_ASAP7_75t_R ID_EX___U353 ( .A(ID_EX__n773), .Y(ID_EX__n266) );
  BUFx2_ASAP7_75t_R ID_EX___U354 ( .A(ID_EX__n780), .Y(ID_EX__n267) );
  BUFx2_ASAP7_75t_R ID_EX___U355 ( .A(ID_EX__n698), .Y(ID_EX__n268) );
  BUFx2_ASAP7_75t_R ID_EX___U356 ( .A(ID_EX__n695), .Y(ID_EX__n269) );
  BUFx2_ASAP7_75t_R ID_EX___U357 ( .A(ID_EX__n688), .Y(ID_EX__n270) );
  BUFx2_ASAP7_75t_R ID_EX___U358 ( .A(ID_EX__n685), .Y(ID_EX__n271) );
  BUFx2_ASAP7_75t_R ID_EX___U359 ( .A(ID_EX__n682), .Y(ID_EX__n272) );
  BUFx2_ASAP7_75t_R ID_EX___U360 ( .A(ID_EX__n669), .Y(ID_EX__n273) );
  BUFx2_ASAP7_75t_R ID_EX___U361 ( .A(ID_EX__n710), .Y(ID_EX__n274) );
  BUFx2_ASAP7_75t_R ID_EX___U362 ( .A(ID_EX__n625), .Y(ID_EX__n275) );
  BUFx2_ASAP7_75t_R ID_EX___U364 ( .A(ID_EX__n631), .Y(ID_EX__n276) );
  BUFx2_ASAP7_75t_R ID_EX___U365 ( .A(ID_EX__n665), .Y(ID_EX__n277) );
  INVx1_ASAP7_75t_R ID_EX___U366 ( .A(ID_EX__n628), .Y(ID_EX__n278) );
  AND2x4_ASAP7_75t_R ID_EX___U367 ( .A(IF_ID_inst[27]), .B(ID_EX__n581), .Y(ID_EX__n694) );
  INVx1_ASAP7_75t_R ID_EX___U368 ( .A(ID_EX__n694), .Y(ID_EX__n279) );
  AND2x4_ASAP7_75t_R ID_EX___U369 ( .A(IF_ID_inst_addr[1]), .B(ID_EX__n574), .Y(ID_EX__n700) );
  INVx1_ASAP7_75t_R ID_EX___U370 ( .A(ID_EX__n700), .Y(ID_EX__n280) );
  AND2x2_ASAP7_75t_R ID_EX___U371 ( .A(IF_ID_inst_addr[21]), .B(ID_EX__n576), .Y(ID_EX__n722) );
  INVx1_ASAP7_75t_R ID_EX___U372 ( .A(ID_EX__n221), .Y(ID_EX__n281) );
  AND2x2_ASAP7_75t_R ID_EX___U373 ( .A(IF_ID_inst_addr[17]), .B(ID_EX__n580), .Y(ID_EX__n718) );
  INVx1_ASAP7_75t_R ID_EX___U374 ( .A(ID_EX__n209), .Y(ID_EX__n282) );
  AND2x2_ASAP7_75t_R ID_EX___U375 ( .A(IF_ID_inst_addr[8]), .B(ID_EX__n614), .Y(ID_EX__n708) );
  INVx1_ASAP7_75t_R ID_EX___U376 ( .A(ID_EX__n207), .Y(ID_EX__n283) );
  AND2x2_ASAP7_75t_R ID_EX___U377 ( .A(IF_ID_inst_addr[4]), .B(ID_EX__n128), .Y(ID_EX__n704) );
  INVx1_ASAP7_75t_R ID_EX___U378 ( .A(ID_EX__n181), .Y(ID_EX__n284) );
  AND2x2_ASAP7_75t_R ID_EX___U379 ( .A(ID_imm[12]), .B(ID_EX__n586), .Y(ID_EX__n645) );
  INVx1_ASAP7_75t_R ID_EX___U380 ( .A(ID_EX__n136), .Y(ID_EX__n285) );
  BUFx6f_ASAP7_75t_R ID_EX___U381 ( .A(ID_EX__n409), .Y(ID_EX_rs1[1]) );
  BUFx2_ASAP7_75t_R ID_EX___U382 ( .A(ID_EX__n768), .Y(ID_EX__n287) );
  BUFx2_ASAP7_75t_R ID_EX___U383 ( .A(ID_EX__n750), .Y(ID_EX__n288) );
  BUFx2_ASAP7_75t_R ID_EX___U384 ( .A(ID_EX__n792), .Y(ID_EX__n289) );
  BUFx2_ASAP7_75t_R ID_EX___U385 ( .A(ID_EX__n741), .Y(ID_EX__n290) );
  BUFx2_ASAP7_75t_R ID_EX___U386 ( .A(ID_EX__n759), .Y(ID_EX__n291) );
  BUFx2_ASAP7_75t_R ID_EX___U387 ( .A(ID_EX__n293), .Y(ID_EX_read_reg_data_2[4]) );
  BUFx2_ASAP7_75t_R ID_EX___U388 ( .A(ID_EX__n799), .Y(ID_EX__n293) );
  BUFx2_ASAP7_75t_R ID_EX___U389 ( .A(ID_EX__n295), .Y(ID_EX_read_reg_data_2[3]) );
  BUFx2_ASAP7_75t_R ID_EX___U390 ( .A(ID_EX__n800), .Y(ID_EX__n295) );
  BUFx3_ASAP7_75t_R ID_EX___U391 ( .A(ID_EX__n297), .Y(ID_EX__n296) );
  BUFx2_ASAP7_75t_R ID_EX___U392 ( .A(ID_EX__n825), .Y(ID_EX__n297) );
  BUFx3_ASAP7_75t_R ID_EX___U393 ( .A(ID_EX__n299), .Y(ID_EX__n298) );
  BUFx2_ASAP7_75t_R ID_EX___U394 ( .A(ID_EX__n827), .Y(ID_EX__n299) );
  BUFx6f_ASAP7_75t_R ID_EX___U395 ( .A(ID_EX__n418), .Y(ID_EX__n300) );
  BUFx3_ASAP7_75t_R ID_EX___U396 ( .A(ID_EX__n302), .Y(ID_EX__n301) );
  BUFx2_ASAP7_75t_R ID_EX___U397 ( .A(ID_EX__n837), .Y(ID_EX__n302) );
  BUFx6f_ASAP7_75t_R ID_EX___U398 ( .A(ID_EX__n472), .Y(ID_EX__n303) );
  BUFx3_ASAP7_75t_R ID_EX___U399 ( .A(ID_EX__n305), .Y(ID_EX__n304) );
  BUFx2_ASAP7_75t_R ID_EX___U400 ( .A(ID_EX__n840), .Y(ID_EX__n305) );
  BUFx6f_ASAP7_75t_R ID_EX___U401 ( .A(ID_EX__n468), .Y(ID_EX__n306) );
  BUFx6f_ASAP7_75t_R ID_EX___U402 ( .A(ID_EX__n413), .Y(ID_EX_inst_12_) );
  AND2x2_ASAP7_75t_R ID_EX___U403 ( .A(n9), .B(ID_EX__n573), .Y(ID_EX__n632) );
  INVx1_ASAP7_75t_R ID_EX___U404 ( .A(ID_EX__n224), .Y(ID_EX__n307) );
  BUFx10_ASAP7_75t_R ID_EX___U405 ( .A(ID_EX__n817), .Y(ID_EX__n411) );
  BUFx6f_ASAP7_75t_R ID_EX___U406 ( .A(ID_EX__n309), .Y(ID_EX_inst_6_) );
  BUFx4f_ASAP7_75t_R ID_EX___U407 ( .A(ID_EX__n188), .Y(ID_EX__n309) );
  BUFx2_ASAP7_75t_R ID_EX___U408 ( .A(ID_EX__n692), .Y(ID_EX__n310) );
  BUFx2_ASAP7_75t_R ID_EX___U409 ( .A(ID_EX__n687), .Y(ID_EX__n311) );
  BUFx2_ASAP7_75t_R ID_EX___U410 ( .A(ID_EX__n635), .Y(ID_EX__n312) );
  AND2x2_ASAP7_75t_R ID_EX___U411 ( .A(ID_EX__n617), .B(ID_MemToReg), .Y(ID_EX__n639) );
  AND2x4_ASAP7_75t_R ID_EX___U412 ( .A(IF_ID_inst[30]), .B(ID_EX__n582), .Y(ID_EX__n697) );
  INVx1_ASAP7_75t_R ID_EX___U413 ( .A(ID_EX__n697), .Y(ID_EX__n314) );
  AND2x4_ASAP7_75t_R ID_EX___U414 ( .A(IF_ID_inst_addr[31]), .B(ID_EX__n579), .Y(ID_EX__n733) );
  INVx1_ASAP7_75t_R ID_EX___U415 ( .A(ID_EX__n733), .Y(ID_EX__n315) );
  AND2x4_ASAP7_75t_R ID_EX___U416 ( .A(IF_ID_inst_addr[26]), .B(ID_EX__n577), .Y(ID_EX__n728) );
  INVx1_ASAP7_75t_R ID_EX___U417 ( .A(ID_EX__n728), .Y(ID_EX__n316) );
  AND2x4_ASAP7_75t_R ID_EX___U418 ( .A(IF_ID_inst_addr[0]), .B(ID_EX__n574), .Y(ID_EX__n699) );
  INVx1_ASAP7_75t_R ID_EX___U419 ( .A(ID_EX__n699), .Y(ID_EX__n317) );
  AND2x2_ASAP7_75t_R ID_EX___U420 ( .A(IF_ID_rd[4]), .B(ID_EX__n95), .Y(ID_EX__n627) );
  INVx1_ASAP7_75t_R ID_EX___U421 ( .A(ID_EX__n223), .Y(ID_EX__n318) );
  AND2x2_ASAP7_75t_R ID_EX___U422 ( .A(IF_ID_rd[1]), .B(ID_EX__n573), .Y(ID_EX__n624) );
  INVx1_ASAP7_75t_R ID_EX___U423 ( .A(ID_EX__n208), .Y(ID_EX__n319) );
  AND2x2_ASAP7_75t_R ID_EX___U424 ( .A(IF_ID_inst_addr[27]), .B(ID_EX__n578), .Y(ID_EX__n729) );
  INVx1_ASAP7_75t_R ID_EX___U425 ( .A(ID_EX__n219), .Y(ID_EX__n320) );
  AND2x2_ASAP7_75t_R ID_EX___U426 ( .A(IF_ID_inst_addr[23]), .B(ID_EX__n576), .Y(ID_EX__n725) );
  INVx1_ASAP7_75t_R ID_EX___U427 ( .A(ID_EX__n180), .Y(ID_EX__n321) );
  AND2x2_ASAP7_75t_R ID_EX___U428 ( .A(IF_ID_inst_addr[12]), .B(ID_EX__n575), .Y(ID_EX__n712) );
  INVx1_ASAP7_75t_R ID_EX___U429 ( .A(ID_EX__n210), .Y(ID_EX__n322) );
  AND2x2_ASAP7_75t_R ID_EX___U430 ( .A(IF_ID_inst_addr[10]), .B(ID_EX__n607), .Y(ID_EX__n710) );
  INVx1_ASAP7_75t_R ID_EX___U431 ( .A(ID_EX__n274), .Y(ID_EX__n323) );
  AND2x2_ASAP7_75t_R ID_EX___U432 ( .A(IF_ID_inst_addr[7]), .B(ID_EX__n605), .Y(ID_EX__n707) );
  INVx1_ASAP7_75t_R ID_EX___U433 ( .A(ID_EX__n250), .Y(ID_EX__n324) );
  AND2x2_ASAP7_75t_R ID_EX___U434 ( .A(n15), .B(ID_EX__n571), .Y(ID_EX__n637) );
  INVx1_ASAP7_75t_R ID_EX___U435 ( .A(ID_EX__n255), .Y(ID_EX__n325) );
  BUFx2_ASAP7_75t_R ID_EX___U436 ( .A(ID_EX__n771), .Y(ID_EX__n326) );
  BUFx2_ASAP7_75t_R ID_EX___U437 ( .A(ID_EX__n767), .Y(ID_EX__n327) );
  BUFx2_ASAP7_75t_R ID_EX___U438 ( .A(ID_EX__n769), .Y(ID_EX__n328) );
  BUFx2_ASAP7_75t_R ID_EX___U439 ( .A(ID_EX__n330), .Y(ID_EX_read_reg_data_1[5]) );
  BUFx2_ASAP7_75t_R ID_EX___U440 ( .A(ID_EX__n766), .Y(ID_EX__n330) );
  BUFx2_ASAP7_75t_R ID_EX___U441 ( .A(ID_EX__n332), .Y(ID_EX_read_reg_data_1[11]) );
  BUFx2_ASAP7_75t_R ID_EX___U442 ( .A(ID_EX__n760), .Y(ID_EX__n332) );
  BUFx2_ASAP7_75t_R ID_EX___U443 ( .A(ID_EX__n747), .Y(ID_EX__n333) );
  BUFx2_ASAP7_75t_R ID_EX___U444 ( .A(ID_EX__n819), .Y(ID_EX__n334) );
  BUFx3_ASAP7_75t_R ID_EX___U445 ( .A(ID_EX__n336), .Y(ID_EX__n335) );
  BUFx2_ASAP7_75t_R ID_EX___U446 ( .A(ID_EX__n826), .Y(ID_EX__n336) );
  AND2x2_ASAP7_75t_R ID_EX___U447 ( .A(ID_EX__n583), .B(ID_imm[1]), .Y(ID_EX__n670) );
  INVx1_ASAP7_75t_R ID_EX___U448 ( .A(ID_EX__n629), .Y(ID_EX__n337) );
  BUFx12f_ASAP7_75t_R ID_EX___U449 ( .A(ID_EX__n806), .Y(ID_EX__n338) );
  BUFx2_ASAP7_75t_R ID_EX___U450 ( .A(ID_EX__n716), .Y(ID_EX__n340) );
  BUFx3_ASAP7_75t_R ID_EX___U451 ( .A(ID_EX__n535), .Y(ID_EX_read_reg_data_1[23]) );
  AND2x2_ASAP7_75t_R ID_EX___U452 ( .A(IF_ID_inst[20]), .B(ID_EX__n615), .Y(ID_EX__n687) );
  INVx1_ASAP7_75t_R ID_EX___U453 ( .A(ID_EX__n311), .Y(ID_EX__n341) );
  AND2x4_ASAP7_75t_R ID_EX___U454 ( .A(IF_ID_inst_addr[30]), .B(ID_EX__n579), .Y(ID_EX__n732) );
  INVx1_ASAP7_75t_R ID_EX___U455 ( .A(ID_EX__n732), .Y(ID_EX__n342) );
  AND2x4_ASAP7_75t_R ID_EX___U456 ( .A(IF_ID_inst_addr[24]), .B(ID_EX__n577), .Y(ID_EX__n726) );
  INVx1_ASAP7_75t_R ID_EX___U457 ( .A(ID_EX__n726), .Y(ID_EX__n343) );
  AND2x4_ASAP7_75t_R ID_EX___U458 ( .A(IF_ID_inst_addr[19]), .B(ID_EX__n570), .Y(ID_EX__n720) );
  INVx1_ASAP7_75t_R ID_EX___U459 ( .A(ID_EX__n720), .Y(ID_EX__n344) );
  AND2x4_ASAP7_75t_R ID_EX___U460 ( .A(IF_ID_inst_addr[2]), .B(ID_EX__n574), .Y(ID_EX__n701) );
  INVx1_ASAP7_75t_R ID_EX___U461 ( .A(ID_EX__n701), .Y(ID_EX__n345) );
  AND2x2_ASAP7_75t_R ID_EX___U462 ( .A(IF_ID_rd[3]), .B(ID_EX__n112), .Y(ID_EX__n626) );
  INVx1_ASAP7_75t_R ID_EX___U463 ( .A(ID_EX__n252), .Y(ID_EX__n346) );
  AND2x2_ASAP7_75t_R ID_EX___U464 ( .A(IF_ID_rd[0]), .B(ID_EX__n115), .Y(ID_EX__n734) );
  INVx1_ASAP7_75t_R ID_EX___U465 ( .A(ID_EX__n253), .Y(ID_EX__n347) );
  AND2x2_ASAP7_75t_R ID_EX___U466 ( .A(IF_ID_inst[31]), .B(ID_EX__n583), .Y(ID_EX__n698) );
  INVx1_ASAP7_75t_R ID_EX___U467 ( .A(ID_EX__n268), .Y(ID_EX__n348) );
  AND2x4_ASAP7_75t_R ID_EX___U468 ( .A(IF_ID_inst[23]), .B(ID_EX__n601), .Y(ID_EX__n690) );
  INVx1_ASAP7_75t_R ID_EX___U469 ( .A(ID_EX__n690), .Y(ID_EX__n349) );
  AND2x4_ASAP7_75t_R ID_EX___U470 ( .A(IF_ID_inst[17]), .B(ID_EX__n599), .Y(ID_EX__n684) );
  INVx1_ASAP7_75t_R ID_EX___U471 ( .A(ID_EX__n684), .Y(ID_EX__n350) );
  AND2x4_ASAP7_75t_R ID_EX___U472 ( .A(IF_ID_inst[11]), .B(ID_EX__n129), .Y(ID_EX__n677) );
  INVx1_ASAP7_75t_R ID_EX___U473 ( .A(ID_EX__n677), .Y(ID_EX__n351) );
  AND2x2_ASAP7_75t_R ID_EX___U474 ( .A(IF_ID_inst_addr[29]), .B(ID_EX__n578), .Y(ID_EX__n731) );
  INVx1_ASAP7_75t_R ID_EX___U475 ( .A(ID_EX__n206), .Y(ID_EX__n352) );
  AND2x2_ASAP7_75t_R ID_EX___U476 ( .A(IF_ID_inst_addr[22]), .B(ID_EX__n576), .Y(ID_EX__n723) );
  INVx1_ASAP7_75t_R ID_EX___U477 ( .A(ID_EX__n170), .Y(ID_EX__n353) );
  BUFx2_ASAP7_75t_R ID_EX___U478 ( .A(ID_EX__n355), .Y(ID_EX_read_reg_data_1[25]) );
  BUFx2_ASAP7_75t_R ID_EX___U479 ( .A(ID_EX__n746), .Y(ID_EX__n355) );
  BUFx2_ASAP7_75t_R ID_EX___U480 ( .A(ID_EX__n753), .Y(ID_EX__n356) );
  BUFx2_ASAP7_75t_R ID_EX___U481 ( .A(ID_EX__n358), .Y(ID_EX_read_reg_data_1[22]) );
  BUFx2_ASAP7_75t_R ID_EX___U482 ( .A(ID_EX__n749), .Y(ID_EX__n358) );
  BUFx2_ASAP7_75t_R ID_EX___U483 ( .A(ID_EX__n758), .Y(ID_EX__n359) );
  BUFx2_ASAP7_75t_R ID_EX___U484 ( .A(ID_EX__n775), .Y(ID_EX__n360) );
  BUFx2_ASAP7_75t_R ID_EX___U485 ( .A(ID_EX__n757), .Y(ID_EX__n362) );
  BUFx2_ASAP7_75t_R ID_EX___U486 ( .A(ID_EX__n743), .Y(ID_EX__n364) );
  BUFx2_ASAP7_75t_R ID_EX___U487 ( .A(ID_EX__n744), .Y(ID_EX__n365) );
  AND2x2_ASAP7_75t_R ID_EX___U488 ( .A(ID_imm[30]), .B(ID_EX__n575), .Y(ID_EX__n663) );
  BUFx2_ASAP7_75t_R ID_EX___U489 ( .A(ID_EX__n367), .Y(ID_EX_read_reg_data_2[26]) );
  BUFx2_ASAP7_75t_R ID_EX___U490 ( .A(ID_EX__n777), .Y(ID_EX__n367) );
  BUFx2_ASAP7_75t_R ID_EX___U491 ( .A(ID_EX__n812), .Y(ID_EX_inst_29_) );
  AND2x2_ASAP7_75t_R ID_EX___U492 ( .A(n7), .B(ID_EX__n594), .Y(ID_EX__n666) );
  INVx1_ASAP7_75t_R ID_EX___U493 ( .A(ID_EX__n247), .Y(ID_EX__n369) );
  AND2x2_ASAP7_75t_R ID_EX___U494 ( .A(n10), .B(ID_EX__n572), .Y(ID_EX__n630) );
  INVx1_ASAP7_75t_R ID_EX___U495 ( .A(ID_EX__n149), .Y(ID_EX__n370) );
  BUFx4f_ASAP7_75t_R ID_EX___U496 ( .A(ID_EX__n372), .Y(ID_EX__n371) );
  BUFx3_ASAP7_75t_R ID_EX___U497 ( .A(ID_EX__n818), .Y(ID_EX__n372) );
  BUFx6f_ASAP7_75t_R ID_EX___U498 ( .A(ID_EX__n371), .Y(ID_EX__n562) );
  BUFx4f_ASAP7_75t_R ID_EX___U499 ( .A(ID_EX__n236), .Y(ID_EX__n374) );
  AND2x2_ASAP7_75t_R ID_EX___U500 ( .A(IF_ID_rd[2]), .B(ID_EX__n111), .Y(ID_EX__n625) );
  INVx1_ASAP7_75t_R ID_EX___U501 ( .A(ID_EX__n275), .Y(ID_EX__n375) );
  AND2x4_ASAP7_75t_R ID_EX___U502 ( .A(IF_ID_inst[22]), .B(ID_EX__n577), .Y(ID_EX__n689) );
  INVx1_ASAP7_75t_R ID_EX___U503 ( .A(ID_EX__n689), .Y(ID_EX__n376) );
  AND2x4_ASAP7_75t_R ID_EX___U504 ( .A(IF_ID_inst[16]), .B(ID_EX__n599), .Y(ID_EX__n683) );
  INVx1_ASAP7_75t_R ID_EX___U505 ( .A(ID_EX__n683), .Y(ID_EX__n377) );
  AND2x4_ASAP7_75t_R ID_EX___U506 ( .A(IF_ID_inst[10]), .B(ID_EX__n608), .Y(ID_EX__n676) );
  INVx1_ASAP7_75t_R ID_EX___U507 ( .A(ID_EX__n676), .Y(ID_EX__n378) );
  AND2x4_ASAP7_75t_R ID_EX___U508 ( .A(IF_ID_inst[8]), .B(ID_EX__n125), .Y(ID_EX__n674) );
  INVx1_ASAP7_75t_R ID_EX___U509 ( .A(ID_EX__n674), .Y(ID_EX__n379) );
  AND2x2_ASAP7_75t_R ID_EX___U510 ( .A(IF_ID_inst_addr[25]), .B(ID_EX__n577), .Y(ID_EX__n727) );
  INVx1_ASAP7_75t_R ID_EX___U511 ( .A(ID_EX__n220), .Y(ID_EX__n380) );
  AND2x2_ASAP7_75t_R ID_EX___U512 ( .A(IF_ID_inst_addr[18]), .B(ID_EX__n128), .Y(ID_EX__n719) );
  INVx1_ASAP7_75t_R ID_EX___U513 ( .A(ID_EX__n173), .Y(ID_EX__n381) );
  AND2x2_ASAP7_75t_R ID_EX___U514 ( .A(IF_ID_inst_addr[15]), .B(ID_EX__n575), .Y(ID_EX__n716) );
  INVx1_ASAP7_75t_R ID_EX___U515 ( .A(ID_EX__n340), .Y(ID_EX__n382) );
  AND2x2_ASAP7_75t_R ID_EX___U516 ( .A(IF_ID_inst_addr[13]), .B(ID_EX__n575), .Y(ID_EX__n714) );
  INVx1_ASAP7_75t_R ID_EX___U517 ( .A(ID_EX__n248), .Y(ID_EX__n383) );
  AND2x2_ASAP7_75t_R ID_EX___U518 ( .A(IF_ID_inst_addr[5]), .B(ID_EX__n158), .Y(ID_EX__n705) );
  INVx1_ASAP7_75t_R ID_EX___U519 ( .A(ID_EX__n251), .Y(ID_EX__n384) );
  AND2x2_ASAP7_75t_R ID_EX___U520 ( .A(IF_ID_inst[6]), .B(ID_EX__n580), .Y(ID_EX__n672) );
  INVx1_ASAP7_75t_R ID_EX___U521 ( .A(ID_EX__n254), .Y(ID_EX__n385) );
  BUFx2_ASAP7_75t_R ID_EX___U522 ( .A(ID_EX__n755), .Y(ID_EX__n386) );
  BUFx2_ASAP7_75t_R ID_EX___U523 ( .A(ID_EX__n765), .Y(ID_EX__n387) );
  BUFx2_ASAP7_75t_R ID_EX___U524 ( .A(ID_EX__n763), .Y(ID_EX__n388) );
  BUFx2_ASAP7_75t_R ID_EX___U525 ( .A(ID_EX__n754), .Y(ID_EX__n389) );
  BUFx2_ASAP7_75t_R ID_EX___U526 ( .A(ID_EX__n762), .Y(ID_EX__n390) );
  BUFx2_ASAP7_75t_R ID_EX___U527 ( .A(ID_EX__n748), .Y(ID_EX__n391) );
  BUFx2_ASAP7_75t_R ID_EX___U528 ( .A(ID_EX__n742), .Y(ID_EX__n392) );
  BUFx2_ASAP7_75t_R ID_EX___U529 ( .A(ID_EX__n801), .Y(ID_EX_read_reg_data_2[2]) );
  BUFx2_ASAP7_75t_R ID_EX___U530 ( .A(ID_EX__n265), .Y(ID_EX_read_reg_data_2[9]) );
  BUFx2_ASAP7_75t_R ID_EX___U531 ( .A(ID_EX__n396), .Y(ID_EX_read_reg_data_2[14]) );
  BUFx2_ASAP7_75t_R ID_EX___U532 ( .A(ID_EX__n789), .Y(ID_EX__n396) );
  BUFx2_ASAP7_75t_R ID_EX___U533 ( .A(ID_EX__n196), .Y(ID_EX_read_reg_data_2[31]) );
  BUFx2_ASAP7_75t_R ID_EX___U534 ( .A(ID_EX__n213), .Y(ID_EX_read_reg_data_2[24]) );
  BUFx2_ASAP7_75t_R ID_EX___U535 ( .A(ID_EX__n400), .Y(ID_EX_read_reg_data_2[19]) );
  BUFx2_ASAP7_75t_R ID_EX___U536 ( .A(ID_EX__n784), .Y(ID_EX__n400) );
  BUFx2_ASAP7_75t_R ID_EX___U537 ( .A(ID_EX__n266), .Y(ID_EX_read_reg_data_2[30]) );
  BUFx2_ASAP7_75t_R ID_EX___U538 ( .A(ID_EX__n403), .Y(ID_EX_read_reg_data_1[18]) );
  BUFx2_ASAP7_75t_R ID_EX___U539 ( .A(ID_EX__n356), .Y(ID_EX__n403) );
  BUFx2_ASAP7_75t_R ID_EX___U540 ( .A(ID_EX__n405), .Y(ID_EX_read_reg_data_1[10]) );
  BUFx2_ASAP7_75t_R ID_EX___U541 ( .A(ID_EX__n264), .Y(ID_EX__n405) );
  AND2x2_ASAP7_75t_R ID_EX___U542 ( .A(IF_ID_inst[0]), .B(ID_EX__n579), .Y(ID_EX__n665) );
  INVx1_ASAP7_75t_R ID_EX___U543 ( .A(ID_EX__n277), .Y(ID_EX__n406) );
  BUFx3_ASAP7_75t_R ID_EX___U544 ( .A(ID_EX__n408), .Y(ID_EX__n407) );
  BUFx2_ASAP7_75t_R ID_EX___U545 ( .A(ID_EX__n838), .Y(ID_EX__n408) );
  BUFx6f_ASAP7_75t_R ID_EX___U546 ( .A(ID_EX__n560), .Y(ID_EX__n409) );
  AND2x2_ASAP7_75t_R ID_EX___U547 ( .A(IF_ID_inst[3]), .B(ID_EX__n613), .Y(ID_EX__n668) );
  INVx1_ASAP7_75t_R ID_EX___U548 ( .A(ID_EX__n169), .Y(ID_EX__n410) );
  BUFx6f_ASAP7_75t_R ID_EX___U549 ( .A(ID_EX__n415), .Y(ID_EX_imm[31]) );
  BUFx4f_ASAP7_75t_R ID_EX___U550 ( .A(ID_EX__n198), .Y(ID_EX__n415) );
  BUFx6f_ASAP7_75t_R ID_EX___U551 ( .A(ID_EX__n417), .Y(ID_EX__n416) );
  BUFx4f_ASAP7_75t_R ID_EX___U552 ( .A(ID_EX__n240), .Y(ID_EX__n417) );
  BUFx6f_ASAP7_75t_R ID_EX___U553 ( .A(ID_EX__n419), .Y(ID_EX__n418) );
  BUFx4f_ASAP7_75t_R ID_EX___U554 ( .A(ID_EX__n298), .Y(ID_EX__n419) );
  BUFx6f_ASAP7_75t_R ID_EX___U555 ( .A(ID_EX__n421), .Y(ID_EX_inst_4_) );
  BUFx4f_ASAP7_75t_R ID_EX___U556 ( .A(ID_EX__n238), .Y(ID_EX__n421) );
  BUFx12f_ASAP7_75t_R ID_EX___U557 ( .A(ID_EX__n423), .Y(ID_EX_imm[30]) );
  BUFx12f_ASAP7_75t_R ID_EX___U558 ( .A(ID_EX__n805), .Y(ID_EX__n423) );
  BUFx12f_ASAP7_75t_R ID_EX___U559 ( .A(ID_EX__n426), .Y(ID_EX_inst_addr[19]) );
  BUFx12f_ASAP7_75t_R ID_EX___U560 ( .A(ID_EX__n832), .Y(ID_EX__n426) );
  BUFx12f_ASAP7_75t_R ID_EX___U561 ( .A(ID_EX__n429), .Y(ID_EX_inst_2_) );
  BUFx12f_ASAP7_75t_R ID_EX___U562 ( .A(ID_EX__n824), .Y(ID_EX__n429) );
  BUFx2_ASAP7_75t_R ID_EX___U563 ( .A(ID_EX__n667), .Y(ID_EX__n430) );
  AND2x4_ASAP7_75t_R ID_EX___U564 ( .A(IF_ID_inst[9]), .B(ID_EX__n126), .Y(ID_EX__n675) );
  INVx1_ASAP7_75t_R ID_EX___U565 ( .A(ID_EX__n675), .Y(ID_EX__n431) );
  AND2x4_ASAP7_75t_R ID_EX___U566 ( .A(IF_ID_inst[7]), .B(ID_EX__n611), .Y(ID_EX__n673) );
  INVx1_ASAP7_75t_R ID_EX___U567 ( .A(ID_EX__n673), .Y(ID_EX__n432) );
  AND2x2_ASAP7_75t_R ID_EX___U568 ( .A(IF_ID_inst[4]), .B(ID_EX__n580), .Y(ID_EX__n669) );
  INVx1_ASAP7_75t_R ID_EX___U569 ( .A(ID_EX__n273), .Y(ID_EX__n433) );
  AND2x2_ASAP7_75t_R ID_EX___U570 ( .A(IF_ID_inst_addr[11]), .B(ID_EX__n140), .Y(ID_EX__n711) );
  INVx1_ASAP7_75t_R ID_EX___U571 ( .A(ID_EX__n249), .Y(ID_EX__n434) );
  BUFx2_ASAP7_75t_R ID_EX___U572 ( .A(ID_EX__n782), .Y(ID_EX_read_reg_data_2[21]) );
  BUFx2_ASAP7_75t_R ID_EX___U573 ( .A(ID_EX__n798), .Y(ID_EX_read_reg_data_2[5]) );
  BUFx2_ASAP7_75t_R ID_EX___U574 ( .A(ID_EX__n751), .Y(ID_EX__n435) );
  BUFx2_ASAP7_75t_R ID_EX___U575 ( .A(ID_EX__n770), .Y(ID_EX__n436) );
  BUFx2_ASAP7_75t_R ID_EX___U576 ( .A(ID_EX__n740), .Y(ID_EX__n437) );
  BUFx2_ASAP7_75t_R ID_EX___U577 ( .A(ID_EX__n764), .Y(ID_EX__n438) );
  BUFx2_ASAP7_75t_R ID_EX___U578 ( .A(ID_EX__n756), .Y(ID_EX__n439) );
  BUFx2_ASAP7_75t_R ID_EX___U579 ( .A(ID_EX__n752), .Y(ID_EX__n440) );
  BUFx2_ASAP7_75t_R ID_EX___U580 ( .A(ID_EX__n786), .Y(ID_EX_read_reg_data_2[17]) );
  BUFx2_ASAP7_75t_R ID_EX___U581 ( .A(ID_EX__n745), .Y(ID_EX__n441) );
  BUFx2_ASAP7_75t_R ID_EX___U582 ( .A(ID_EX__n186), .Y(ID_EX_read_reg_data_2[18]) );
  BUFx2_ASAP7_75t_R ID_EX___U583 ( .A(ID_EX__n233), .Y(ID_EX_read_reg_data_2[1]) );
  BUFx2_ASAP7_75t_R ID_EX___U584 ( .A(ID_EX__n289), .Y(ID_EX_read_reg_data_2[11]) );
  BUFx2_ASAP7_75t_R ID_EX___U585 ( .A(ID_EX__n212), .Y(ID_EX_read_reg_data_2[13]) );
  BUFx2_ASAP7_75t_R ID_EX___U586 ( .A(ID_EX__n360), .Y(ID_EX_read_reg_data_2[28]) );
  BUFx2_ASAP7_75t_R ID_EX___U587 ( .A(ID_EX__n788), .Y(ID_EX_read_reg_data_2[15]) );
  BUFx2_ASAP7_75t_R ID_EX___U588 ( .A(ID_EX__n267), .Y(ID_EX_read_reg_data_2[23]) );
  BUFx2_ASAP7_75t_R ID_EX___U589 ( .A(ID_EX__n813), .Y(ID_EX_inst_28_) );
  BUFx2_ASAP7_75t_R ID_EX___U590 ( .A(ID_EX__n451), .Y(ID_EX_MemWrite) );
  BUFx2_ASAP7_75t_R ID_EX___U591 ( .A(ID_EX__n737), .Y(ID_EX__n451) );
  BUFx2_ASAP7_75t_R ID_EX___U592 ( .A(ID_EX__n453), .Y(ID_EX_read_reg_data_1[21]) );
  BUFx2_ASAP7_75t_R ID_EX___U593 ( .A(ID_EX__n288), .Y(ID_EX__n453) );
  BUFx2_ASAP7_75t_R ID_EX___U594 ( .A(ID_EX__n455), .Y(ID_EX_read_reg_data_1[13]) );
  BUFx2_ASAP7_75t_R ID_EX___U595 ( .A(ID_EX__n359), .Y(ID_EX__n455) );
  BUFx2_ASAP7_75t_R ID_EX___U596 ( .A(ID_EX__n457), .Y(ID_EX_read_reg_data_1[17]) );
  BUFx2_ASAP7_75t_R ID_EX___U597 ( .A(ID_EX__n389), .Y(ID_EX__n457) );
  BUFx2_ASAP7_75t_R ID_EX___U598 ( .A(ID_EX__n459), .Y(ID_EX_read_reg_data_1[29]) );
  BUFx2_ASAP7_75t_R ID_EX___U599 ( .A(ID_EX__n392), .Y(ID_EX__n459) );
  AND2x2_ASAP7_75t_R ID_EX___U600 ( .A(IF_ID_inst[29]), .B(ID_EX__n582), .Y(ID_EX__n696) );
  INVx1_ASAP7_75t_R ID_EX___U601 ( .A(ID_EX__n244), .Y(ID_EX__n460) );
  AND2x2_ASAP7_75t_R ID_EX___U602 ( .A(IF_ID_inst[26]), .B(ID_EX__n581), .Y(ID_EX__n693) );
  INVx1_ASAP7_75t_R ID_EX___U603 ( .A(ID_EX__n245), .Y(ID_EX__n461) );
  AND2x2_ASAP7_75t_R ID_EX___U604 ( .A(IF_ID_inst[19]), .B(ID_EX__n599), .Y(ID_EX__n686) );
  INVx1_ASAP7_75t_R ID_EX___U605 ( .A(ID_EX__n246), .Y(ID_EX__n462) );
  BUFx3_ASAP7_75t_R ID_EX___U606 ( .A(ID_EX__n464), .Y(ID_EX__n463) );
  BUFx2_ASAP7_75t_R ID_EX___U607 ( .A(ID_EX__n839), .Y(ID_EX__n464) );
  BUFx6f_ASAP7_75t_R ID_EX___U608 ( .A(ID_EX__n558), .Y(ID_EX_rs1[0]) );
  INVx1_ASAP7_75t_R ID_EX___U609 ( .A(ID_EX__n633), .Y(ID_EX__n466) );
  AND2x2_ASAP7_75t_R ID_EX___U610 ( .A(IF_ID_rs1[3]), .B(ID_EX__n572), .Y(ID_EX__n631) );
  INVx1_ASAP7_75t_R ID_EX___U611 ( .A(ID_EX__n276), .Y(ID_EX__n467) );
  BUFx6f_ASAP7_75t_R ID_EX___U612 ( .A(ID_EX__n469), .Y(ID_EX__n468) );
  BUFx4f_ASAP7_75t_R ID_EX___U613 ( .A(ID_EX__n304), .Y(ID_EX__n469) );
  BUFx6f_ASAP7_75t_R ID_EX___U614 ( .A(ID_EX__n471), .Y(ID_EX__n470) );
  BUFx4f_ASAP7_75t_R ID_EX___U615 ( .A(ID_EX__n214), .Y(ID_EX__n471) );
  BUFx6f_ASAP7_75t_R ID_EX___U616 ( .A(ID_EX__n473), .Y(ID_EX__n472) );
  BUFx4f_ASAP7_75t_R ID_EX___U617 ( .A(ID_EX__n301), .Y(ID_EX__n473) );
  BUFx6f_ASAP7_75t_R ID_EX___U618 ( .A(ID_EX__n475), .Y(ID_EX_inst_5_) );
  BUFx4f_ASAP7_75t_R ID_EX___U619 ( .A(ID_EX__n200), .Y(ID_EX__n475) );
  BUFx12f_ASAP7_75t_R ID_EX___U620 ( .A(ID_EX__n483), .Y(ID_EX_imm[29]) );
  BUFx12f_ASAP7_75t_R ID_EX___U621 ( .A(ID_EX__n338), .Y(ID_EX__n483) );
  BUFx2_ASAP7_75t_R ID_EX___U622 ( .A(ID_EX__n778), .Y(ID_EX_read_reg_data_2[25]) );
  BUFx2_ASAP7_75t_R ID_EX___U623 ( .A(ID_EX__n781), .Y(ID_EX_read_reg_data_2[22]) );
  BUFx2_ASAP7_75t_R ID_EX___U624 ( .A(ID_EX__n783), .Y(ID_EX_read_reg_data_2[20]) );
  BUFx2_ASAP7_75t_R ID_EX___U625 ( .A(ID_EX__n787), .Y(ID_EX_read_reg_data_2[16]) );
  BUFx2_ASAP7_75t_R ID_EX___U626 ( .A(ID_EX__n795), .Y(ID_EX_read_reg_data_2[8]) );
  BUFx2_ASAP7_75t_R ID_EX___U627 ( .A(ID_EX__n797), .Y(ID_EX_read_reg_data_2[6]) );
  BUFx2_ASAP7_75t_R ID_EX___U628 ( .A(ID_EX__n803), .Y(ID_EX_read_reg_data_2[0]) );
  BUFx2_ASAP7_75t_R ID_EX___U629 ( .A(ID_EX__n793), .Y(ID_EX_read_reg_data_2[10]) );
  BUFx2_ASAP7_75t_R ID_EX___U630 ( .A(ID_EX__n796), .Y(ID_EX_read_reg_data_2[7]) );
  BUFx2_ASAP7_75t_R ID_EX___U631 ( .A(ID_EX__n776), .Y(ID_EX_read_reg_data_2[27]) );
  BUFx2_ASAP7_75t_R ID_EX___U632 ( .A(ID_EX__n774), .Y(ID_EX_read_reg_data_2[29]) );
  BUFx2_ASAP7_75t_R ID_EX___U633 ( .A(ID_EX__n791), .Y(ID_EX_read_reg_data_2[12]) );
  BUFx2_ASAP7_75t_R ID_EX___U634 ( .A(ID_EX__n501), .Y(ID_EX_MemToReg) );
  BUFx2_ASAP7_75t_R ID_EX___U635 ( .A(ID_EX__n736), .Y(ID_EX__n501) );
  BUFx2_ASAP7_75t_R ID_EX___U636 ( .A(ID_EX__n503), .Y(ID_EX_read_reg_data_1[0]) );
  BUFx2_ASAP7_75t_R ID_EX___U637 ( .A(ID_EX__n326), .Y(ID_EX__n503) );
  BUFx2_ASAP7_75t_R ID_EX___U638 ( .A(ID_EX__n505), .Y(ID_EX_read_reg_data_1[16]) );
  BUFx2_ASAP7_75t_R ID_EX___U639 ( .A(ID_EX__n386), .Y(ID_EX__n505) );
  BUFx2_ASAP7_75t_R ID_EX___U640 ( .A(ID_EX__n507), .Y(ID_EX_read_reg_data_1[6]) );
  BUFx2_ASAP7_75t_R ID_EX___U641 ( .A(ID_EX__n387), .Y(ID_EX__n507) );
  BUFx2_ASAP7_75t_R ID_EX___U642 ( .A(ID_EX__n509), .Y(ID_EX_read_reg_data_1[8]) );
  BUFx2_ASAP7_75t_R ID_EX___U643 ( .A(ID_EX__n388), .Y(ID_EX__n509) );
  BUFx2_ASAP7_75t_R ID_EX___U644 ( .A(ID_EX__n511), .Y(ID_EX_read_reg_data_1[3]) );
  BUFx2_ASAP7_75t_R ID_EX___U645 ( .A(ID_EX__n287), .Y(ID_EX__n511) );
  BUFx2_ASAP7_75t_R ID_EX___U646 ( .A(ID_EX__n513), .Y(ID_EX_read_reg_data_1[20]) );
  BUFx2_ASAP7_75t_R ID_EX___U647 ( .A(ID_EX__n435), .Y(ID_EX__n513) );
  BUFx2_ASAP7_75t_R ID_EX___U648 ( .A(ID_EX__n515), .Y(ID_EX_read_reg_data_1[4]) );
  BUFx2_ASAP7_75t_R ID_EX___U649 ( .A(ID_EX__n327), .Y(ID_EX__n515) );
  BUFx2_ASAP7_75t_R ID_EX___U650 ( .A(ID_EX__n517), .Y(ID_EX_read_reg_data_1[2]) );
  BUFx2_ASAP7_75t_R ID_EX___U651 ( .A(ID_EX__n328), .Y(ID_EX__n517) );
  BUFx2_ASAP7_75t_R ID_EX___U652 ( .A(ID_EX__n519), .Y(ID_EX_read_reg_data_1[1]) );
  BUFx2_ASAP7_75t_R ID_EX___U653 ( .A(ID_EX__n436), .Y(ID_EX__n519) );
  BUFx2_ASAP7_75t_R ID_EX___U654 ( .A(ID_EX__n521), .Y(ID_EX_read_reg_data_1[9]) );
  BUFx2_ASAP7_75t_R ID_EX___U655 ( .A(ID_EX__n390), .Y(ID_EX__n521) );
  BUFx2_ASAP7_75t_R ID_EX___U656 ( .A(ID_EX__n523), .Y(ID_EX_read_reg_data_1[30]) );
  BUFx2_ASAP7_75t_R ID_EX___U657 ( .A(ID_EX__n290), .Y(ID_EX__n523) );
  BUFx2_ASAP7_75t_R ID_EX___U658 ( .A(ID_EX__n525), .Y(ID_EX_read_reg_data_1[31]) );
  BUFx2_ASAP7_75t_R ID_EX___U659 ( .A(ID_EX__n437), .Y(ID_EX__n525) );
  BUFx2_ASAP7_75t_R ID_EX___U660 ( .A(ID_EX__n527), .Y(ID_EX_read_reg_data_1[7]) );
  BUFx2_ASAP7_75t_R ID_EX___U661 ( .A(ID_EX__n438), .Y(ID_EX__n527) );
  BUFx2_ASAP7_75t_R ID_EX___U662 ( .A(ID_EX__n529), .Y(ID_EX_read_reg_data_1[24]) );
  BUFx2_ASAP7_75t_R ID_EX___U663 ( .A(ID_EX__n333), .Y(ID_EX__n529) );
  BUFx2_ASAP7_75t_R ID_EX___U664 ( .A(ID_EX__n531), .Y(ID_EX_read_reg_data_1[15]) );
  BUFx2_ASAP7_75t_R ID_EX___U665 ( .A(ID_EX__n439), .Y(ID_EX__n531) );
  BUFx2_ASAP7_75t_R ID_EX___U666 ( .A(ID_EX__n533), .Y(ID_EX_read_reg_data_1[19]) );
  BUFx2_ASAP7_75t_R ID_EX___U667 ( .A(ID_EX__n440), .Y(ID_EX__n533) );
  BUFx2_ASAP7_75t_R ID_EX___U668 ( .A(ID_EX__n391), .Y(ID_EX__n535) );
  BUFx2_ASAP7_75t_R ID_EX___U669 ( .A(ID_EX__n537), .Y(ID_EX_read_reg_data_1[12]) );
  BUFx2_ASAP7_75t_R ID_EX___U670 ( .A(ID_EX__n291), .Y(ID_EX__n537) );
  BUFx2_ASAP7_75t_R ID_EX___U671 ( .A(ID_EX__n539), .Y(ID_EX_read_reg_data_1[14]) );
  BUFx2_ASAP7_75t_R ID_EX___U672 ( .A(ID_EX__n362), .Y(ID_EX__n539) );
  BUFx2_ASAP7_75t_R ID_EX___U673 ( .A(ID_EX__n541), .Y(ID_EX_read_reg_data_1[28]) );
  BUFx2_ASAP7_75t_R ID_EX___U674 ( .A(ID_EX__n364), .Y(ID_EX__n541) );
  BUFx2_ASAP7_75t_R ID_EX___U675 ( .A(ID_EX__n543), .Y(ID_EX_read_reg_data_1[26]) );
  BUFx2_ASAP7_75t_R ID_EX___U676 ( .A(ID_EX__n441), .Y(ID_EX__n543) );
  BUFx2_ASAP7_75t_R ID_EX___U677 ( .A(ID_EX__n545), .Y(ID_EX_read_reg_data_1[27]) );
  BUFx2_ASAP7_75t_R ID_EX___U678 ( .A(ID_EX__n365), .Y(ID_EX__n545) );
  AND2x2_ASAP7_75t_R ID_EX___U679 ( .A(IF_ID_inst[28]), .B(ID_EX__n582), .Y(ID_EX__n695) );
  INVx1_ASAP7_75t_R ID_EX___U680 ( .A(ID_EX__n269), .Y(ID_EX__n546) );
  AND2x2_ASAP7_75t_R ID_EX___U681 ( .A(IF_ID_inst[25]), .B(ID_EX__n581), .Y(ID_EX__n692) );
  INVx1_ASAP7_75t_R ID_EX___U682 ( .A(ID_EX__n310), .Y(ID_EX__n547) );
  AND2x2_ASAP7_75t_R ID_EX___U683 ( .A(IF_ID_inst[21]), .B(ID_EX__n579), .Y(ID_EX__n688) );
  INVx1_ASAP7_75t_R ID_EX___U684 ( .A(ID_EX__n270), .Y(ID_EX__n548) );
  AND2x2_ASAP7_75t_R ID_EX___U685 ( .A(IF_ID_inst[12]), .B(ID_EX__n572), .Y(ID_EX__n678) );
  INVx1_ASAP7_75t_R ID_EX___U686 ( .A(ID_EX__n204), .Y(ID_EX__n549) );
  AND2x2_ASAP7_75t_R ID_EX___U687 ( .A(IF_ID_inst[18]), .B(ID_EX__n587), .Y(ID_EX__n685) );
  INVx1_ASAP7_75t_R ID_EX___U688 ( .A(ID_EX__n271), .Y(ID_EX__n550) );
  AND2x2_ASAP7_75t_R ID_EX___U689 ( .A(IF_ID_inst[15]), .B(ID_EX__n599), .Y(ID_EX__n682) );
  INVx1_ASAP7_75t_R ID_EX___U690 ( .A(ID_EX__n272), .Y(ID_EX__n551) );
  AND2x2_ASAP7_75t_R ID_EX___U691 ( .A(IF_ID_inst[2]), .B(ID_EX__n583), .Y(ID_EX__n667) );
  INVx1_ASAP7_75t_R ID_EX___U692 ( .A(ID_EX__n430), .Y(ID_EX__n552) );
  BUFx6f_ASAP7_75t_R ID_EX___U693 ( .A(ID_EX__n554), .Y(ID_EX_inst_1_) );
  BUFx4f_ASAP7_75t_R ID_EX___U694 ( .A(ID_EX__n296), .Y(ID_EX__n554) );
  BUFx6f_ASAP7_75t_R ID_EX___U695 ( .A(ID_EX__n556), .Y(ID_EX_inst_0_) );
  BUFx4f_ASAP7_75t_R ID_EX___U696 ( .A(ID_EX__n335), .Y(ID_EX__n556) );
  AND2x2_ASAP7_75t_R ID_EX___U697 ( .A(n44), .B(ID_EX__n570), .Y(ID_EX__n635) );
  INVx1_ASAP7_75t_R ID_EX___U698 ( .A(ID_EX__n312), .Y(ID_EX__n557) );
  BUFx6f_ASAP7_75t_R ID_EX___U699 ( .A(ID_EX__n559), .Y(ID_EX__n558) );
  BUFx4f_ASAP7_75t_R ID_EX___U700 ( .A(ID_EX__n463), .Y(ID_EX__n559) );
  BUFx6f_ASAP7_75t_R ID_EX___U701 ( .A(ID_EX__n561), .Y(ID_EX__n560) );
  BUFx4f_ASAP7_75t_R ID_EX___U702 ( .A(ID_EX__n407), .Y(ID_EX__n561) );
  BUFx12f_ASAP7_75t_R ID_EX___U703 ( .A(ID_EX__n564), .Y(ID_EX_inst_30_) );
  BUFx12f_ASAP7_75t_R ID_EX___U704 ( .A(ID_EX__n243), .Y(ID_EX__n564) );
  BUFx12f_ASAP7_75t_R ID_EX___U705 ( .A(ID_EX__n566), .Y(ID_EX_inst_addr[29]) );
  BUFx12f_ASAP7_75t_R ID_EX___U706 ( .A(ID_EX__n829), .Y(ID_EX__n566) );
  BUFx12f_ASAP7_75t_R ID_EX___U707 ( .A(ID_EX__n568), .Y(ID_EX_inst_addr[30]) );
  BUFx12f_ASAP7_75t_R ID_EX___U708 ( .A(ID_EX__n828), .Y(ID_EX__n568) );
  BUFx12f_ASAP7_75t_R ID_EX___U709 ( .A(ID_EX__n585), .Y(ID_EX__n571) );
  BUFx12f_ASAP7_75t_R ID_EX___U710 ( .A(ID_EX__n592), .Y(ID_EX__n572) );
  BUFx12f_ASAP7_75t_R ID_EX___U711 ( .A(ID_EX__n586), .Y(ID_EX__n573) );
  BUFx12f_ASAP7_75t_R ID_EX___U712 ( .A(ID_EX__n596), .Y(ID_EX__n574) );
  BUFx12f_ASAP7_75t_R ID_EX___U713 ( .A(ID_EX__n612), .Y(ID_EX__n575) );
  BUFx12f_ASAP7_75t_R ID_EX___U714 ( .A(ID_EX__n593), .Y(ID_EX__n576) );
  BUFx12f_ASAP7_75t_R ID_EX___U715 ( .A(ID_EX__n590), .Y(ID_EX__n577) );
  BUFx12f_ASAP7_75t_R ID_EX___U716 ( .A(ID_EX__n591), .Y(ID_EX__n578) );
  BUFx12f_ASAP7_75t_R ID_EX___U717 ( .A(ID_EX__n589), .Y(ID_EX__n579) );
  BUFx12f_ASAP7_75t_R ID_EX___U718 ( .A(ID_EX__n611), .Y(ID_EX__n580) );
  BUFx12f_ASAP7_75t_R ID_EX___U719 ( .A(ID_EX__n588), .Y(ID_EX__n581) );
  BUFx12f_ASAP7_75t_R ID_EX___U720 ( .A(ID_EX__n598), .Y(ID_EX__n582) );
  BUFx12f_ASAP7_75t_R ID_EX___U721 ( .A(ID_EX__n573), .Y(ID_EX__n583) );
  BUFx12f_ASAP7_75t_R ID_EX___U722 ( .A(ID_EX__n604), .Y(ID_EX__n587) );
  BUFx12f_ASAP7_75t_R ID_EX___U723 ( .A(ID_EX__n610), .Y(ID_EX__n588) );
  BUFx12f_ASAP7_75t_R ID_EX___U724 ( .A(ID_EX__n609), .Y(ID_EX__n589) );
  BUFx12f_ASAP7_75t_R ID_EX___U725 ( .A(ID_EX__n157), .Y(ID_EX__n590) );
  BUFx12f_ASAP7_75t_R ID_EX___U726 ( .A(ID_EX__n158), .Y(ID_EX__n591) );
  BUFx12f_ASAP7_75t_R ID_EX___U727 ( .A(ID_EX__n607), .Y(ID_EX__n592) );
  BUFx12f_ASAP7_75t_R ID_EX___U728 ( .A(ID_EX__n606), .Y(ID_EX__n593) );
  BUFx12f_ASAP7_75t_R ID_EX___U729 ( .A(ID_EX__n605), .Y(ID_EX__n594) );
  BUFx12f_ASAP7_75t_R ID_EX___U730 ( .A(ID_EX__n138), .Y(ID_EX__n595) );
  BUFx12f_ASAP7_75t_R ID_EX___U731 ( .A(ID_EX__n139), .Y(ID_EX__n596) );
  BUFx12f_ASAP7_75t_R ID_EX___U732 ( .A(ID_EX__n603), .Y(ID_EX__n597) );
  BUFx12f_ASAP7_75t_R ID_EX___U733 ( .A(ID_EX__n597), .Y(ID_EX__n598) );
  BUFx12f_ASAP7_75t_R ID_EX___U734 ( .A(ID_EX__n602), .Y(ID_EX__n599) );
  BUFx12f_ASAP7_75t_R ID_EX___U735 ( .A(ID_EX__n601), .Y(ID_EX__n600) );      
  OR2x2_ASAP7_75t_R EX___U233 ( .A(ForwardA[0]), .B(EX__n1578), .Y(EX__n140) );


  OAI31xp33_ASAP7_75t_R ALU___U123 ( .A1(ALU__n1373), .A2(ALU__n1400), .A3(ALU__n1401), .B(ALU__n1506), 
        .Y(ALU_zero) );
  OR5x1_ASAP7_75t_R ALU___U124 ( .A(EX_ALU_result[10]), .B(EX_ALU_result[0]), .C(
        EX_ALU_result[12]), .D(EX_ALU_result[11]), .E(ALU__n972), .Y(ALU__n119) );
  OR4x1_ASAP7_75t_R ALU___U125 ( .A(EX_ALU_result[14]), .B(EX_ALU_result[13]), .C(
        EX_ALU_result[16]), .D(EX_ALU_result[15]), .Y(ALU__n120) );
  OR5x1_ASAP7_75t_R ALU___U126 ( .A(EX_ALU_result[18]), .B(EX_ALU_result[17]), .C(
        EX_ALU_result[1]), .D(EX_ALU_result[19]), .E(ALU__n911), .Y(ALU__n118) );
  OR4x1_ASAP7_75t_R ALU___U127 ( .A(EX_ALU_result[21]), .B(EX_ALU_result[20]), .C(
        EX_ALU_result[23]), .D(EX_ALU_result[22]), .Y(ALU__n121) );
  OR3x1_ASAP7_75t_R ALU___U128 ( .A(ALU__n1190), .B(ALU__n1192), .C(ALU__n1191), .Y(ALU__N387) );
  AO22x1_ASAP7_75t_R ALU___U131 ( .A1(ALU__N322), .A2(ALU__n1519), .B1(ALU__N354), .B2(ALU__n1504), .Y(
        n127) );
  OA221x2_ASAP7_75t_R ALU___U134 ( .A1(ALU__n1445), .A2(ALU__n1775), .B1(ALU__n1479), .B2(
        n1091), .C(ALU__n1588), .Y(ALU__n136) );
  OR3x1_ASAP7_75t_R ALU___U135 ( .A(ALU__n993), .B(ALU__n994), .C(ALU__n992), .Y(ALU__N386) );
  OA22x2_ASAP7_75t_R ALU___U140 ( .A1(ALU__n1198), .A2(ALU__n1481), .B1(ALU__n1454), .B2(
        n1010), .Y(ALU__n146) );
  OA221x2_ASAP7_75t_R ALU___U141 ( .A1(ALU__n1198), .A2(ALU__n1432), .B1(ALU__n1470), .B2(
        n1010), .C(ALU__n1594), .Y(ALU__n145) );
  OR3x1_ASAP7_75t_R ALU___U142 ( .A(ALU__n1027), .B(ALU__n1029), .C(ALU__n1028), .Y(ALU__N385) );
  OA22x2_ASAP7_75t_R ALU___U147 ( .A1(ALU__n1358), .A2(ALU__n1480), .B1(ALU__n1454), .B2(
        n1215), .Y(ALU__n152) );
  OA221x2_ASAP7_75t_R ALU___U148 ( .A1(ALU__n1358), .A2(ALU__n1432), .B1(ALU__n1470), .B2(
        n1215), .C(ALU__n1589), .Y(ALU__n151) );
  OR3x1_ASAP7_75t_R ALU___U149 ( .A(ALU__n1228), .B(ALU__n1229), .C(ALU__n1227), .Y(ALU__N384) );
  OA22x2_ASAP7_75t_R ALU___U154 ( .A1(ALU__n1420), .A2(ALU__n1480), .B1(ALU__n1455), .B2(
        n920), .Y(ALU__n158) );
  OA221x2_ASAP7_75t_R ALU___U155 ( .A1(ALU__n1420), .A2(ALU__n1433), .B1(ALU__n1473), .B2(
        n920), .C(ALU__n1591), .Y(ALU__n157) );
  OR3x1_ASAP7_75t_R ALU___U156 ( .A(ALU__n812), .B(ALU__n813), .C(ALU__n811), .Y(ALU__N383) );
  OA22x2_ASAP7_75t_R ALU___U161 ( .A1(ALU__n1362), .A2(ALU__n1482), .B1(ALU__n1455), .B2(
        n1160), .Y(ALU__n164) );
  OA221x2_ASAP7_75t_R ALU___U162 ( .A1(ALU__n1362), .A2(ALU__n1433), .B1(ALU__n1472), .B2(
        n1160), .C(ALU__n1590), .Y(ALU__n163) );
  OR3x1_ASAP7_75t_R ALU___U163 ( .A(ALU__n1231), .B(ALU__n1233), .C(ALU__n1232), .Y(ALU__N382) );
  AO22x1_ASAP7_75t_R ALU___U166 ( .A1(ALU__N317), .A2(ALU__n1518), .B1(ALU__N349), .B2(ALU__n1505), .Y(
        n166) );
  OA22x2_ASAP7_75t_R ALU___U168 ( .A1(ALU__n1419), .A2(ALU__n1480), .B1(ALU__n1455), .B2(
        n1100), .Y(ALU__n170) );
  OA221x2_ASAP7_75t_R ALU___U169 ( .A1(ALU__n1419), .A2(ALU__n1434), .B1(ALU__n1474), .B2(
        n1100), .C(ALU__n1601), .Y(ALU__n169) );
  OR3x1_ASAP7_75t_R ALU___U170 ( .A(ALU__n1086), .B(ALU__n1088), .C(ALU__n1087), .Y(ALU__N381) );
  AO22x1_ASAP7_75t_R ALU___U173 ( .A1(ALU__N316), .A2(ALU__n1518), .B1(ALU__N348), .B2(ALU__n1505), .Y(
        n172) );
  OA22x2_ASAP7_75t_R ALU___U175 ( .A1(ALU__n1385), .A2(ALU__n1481), .B1(ALU__n1456), .B2(ALU__n934), .Y(
        n176) );
  OA221x2_ASAP7_75t_R ALU___U176 ( .A1(ALU__n1385), .A2(ALU__n1434), .B1(ALU__n696), .B2(ALU__n786), .C(
        n379), .Y(ALU__n175) );
  OR3x1_ASAP7_75t_R ALU___U177 ( .A(ALU__n1178), .B(ALU__n1180), .C(ALU__n1179), .Y(ALU__N380) );
  AO22x1_ASAP7_75t_R ALU___U180 ( .A1(ALU__N315), .A2(ALU__n1518), .B1(ALU__N347), .B2(ALU__n1505), .Y(
        n178) );
  OA22x2_ASAP7_75t_R ALU___U182 ( .A1(ALU__n1392), .A2(ALU__n1482), .B1(ALU__n1456), .B2(
        n1064), .Y(ALU__n182) );
  OA221x2_ASAP7_75t_R ALU___U183 ( .A1(ALU__n1392), .A2(ALU__n1435), .B1(ALU__n11), .B2(
        n1064), .C(ALU__n1594), .Y(ALU__n181) );
  OR3x1_ASAP7_75t_R ALU___U184 ( .A(ALU__n1134), .B(ALU__n1136), .C(ALU__n1135), .Y(ALU__N379) );
  OA22x2_ASAP7_75t_R ALU___U189 ( .A1(ALU__n1359), .A2(ALU__n1481), .B1(ALU__n1456), .B2(
        n1178), .Y(ALU__n188) );
  OA221x2_ASAP7_75t_R ALU___U190 ( .A1(ALU__n1359), .A2(ALU__n1437), .B1(ALU__n21), .B2(
        n1178), .C(ALU__n1596), .Y(ALU__n187) );
  OR3x1_ASAP7_75t_R ALU___U191 ( .A(ALU__n1260), .B(ALU__n1262), .C(ALU__n1261), .Y(ALU__N378) );
  AO22x1_ASAP7_75t_R ALU___U194 ( .A1(ALU__N313), .A2(ALU__n1518), .B1(ALU__N345), .B2(ALU__n1505), .Y(
        n190) );
  OA22x2_ASAP7_75t_R ALU___U196 ( .A1(ALU__n1393), .A2(ALU__n1482), .B1(ALU__n1457), .B2(
        n1024), .Y(ALU__n194) );
  OA221x2_ASAP7_75t_R ALU___U197 ( .A1(ALU__n1393), .A2(ALU__n1435), .B1(ALU__n1478), .B2(
        n1024), .C(ALU__n1587), .Y(ALU__n193) );
  OR3x1_ASAP7_75t_R ALU___U198 ( .A(ALU__n836), .B(ALU__n835), .C(ALU__n834), .Y(ALU__N377) );
  OA22x2_ASAP7_75t_R ALU___U203 ( .A1(ALU__n1335), .A2(ALU__n1483), .B1(ALU__n1457), .B2(
        n1225), .Y(ALU__n200) );
  OA221x2_ASAP7_75t_R ALU___U204 ( .A1(ALU__n1335), .A2(ALU__n1436), .B1(ALU__n1479), .B2(
        n1225), .C(ALU__n1594), .Y(ALU__n199) );
  OR3x1_ASAP7_75t_R ALU___U205 ( .A(ALU__n1113), .B(ALU__n1115), .C(ALU__n1114), .Y(ALU__N376) );
  AO22x1_ASAP7_75t_R ALU___U208 ( .A1(ALU__N311), .A2(ALU__n1517), .B1(ALU__N343), .B2(ALU__n1503), .Y(
        n202) );
  OA22x2_ASAP7_75t_R ALU___U210 ( .A1(ALU__n1418), .A2(ALU__n1483), .B1(ALU__n1457), .B2(
        n1068), .Y(ALU__n206) );
  OA221x2_ASAP7_75t_R ALU___U211 ( .A1(ALU__n1418), .A2(ALU__n1436), .B1(ALU__n19), .B2(
        n1068), .C(ALU__n1605), .Y(ALU__n205) );
  OR3x1_ASAP7_75t_R ALU___U212 ( .A(ALU__n896), .B(ALU__n897), .C(ALU__n895), .Y(ALU__N375) );
  OA22x2_ASAP7_75t_R ALU___U217 ( .A1(ALU__n1394), .A2(ALU__n1484), .B1(ALU__n1458), .B2(ALU__n1035), 
        .Y(ALU__n212) );
  OA221x2_ASAP7_75t_R ALU___U218 ( .A1(ALU__n1394), .A2(ALU__n1443), .B1(ALU__n1479), .B2(ALU__n1037), 
        .C(ALU__n1596), .Y(ALU__n211) );
  OR3x1_ASAP7_75t_R ALU___U219 ( .A(ALU__n998), .B(ALU__n997), .C(ALU__n996), .Y(ALU__N374) );
  OA22x2_ASAP7_75t_R ALU___U224 ( .A1(ALU__n1361), .A2(ALU__n1484), .B1(ALU__n1458), .B2(
        n1182), .Y(ALU__n218) );
  OA221x2_ASAP7_75t_R ALU___U225 ( .A1(ALU__n1361), .A2(ALU__n1442), .B1(ALU__n1478), .B2(
        n1182), .C(ALU__n1592), .Y(ALU__n217) );
  OR3x1_ASAP7_75t_R ALU___U226 ( .A(ALU__n1092), .B(ALU__n1091), .C(ALU__n1090), .Y(ALU__N373) );
  OA22x2_ASAP7_75t_R ALU___U231 ( .A1(ALU__n1388), .A2(ALU__n1484), .B1(ALU__n1458), .B2(ALU__n966), .Y(
        n224) );
  OA221x2_ASAP7_75t_R ALU___U232 ( .A1(ALU__n1388), .A2(ALU__n1434), .B1(ALU__n1476), .B2(ALU__n965), 
        .C(ALU__n1595), .Y(ALU__n223) );
  OR3x1_ASAP7_75t_R ALU___U233 ( .A(ALU__n1265), .B(ALU__n1266), .C(ALU__n1264), .Y(ALU__N372) );
  OA22x2_ASAP7_75t_R ALU___U238 ( .A1(ALU__n981), .A2(ALU__n1485), .B1(ALU__n753), .B2(
        n1073), .Y(ALU__n230) );
  OA221x2_ASAP7_75t_R ALU___U239 ( .A1(ALU__n981), .A2(ALU__n1433), .B1(ALU__n1489), .B2(
        n1073), .C(ALU__n1595), .Y(ALU__n229) );
  OR3x1_ASAP7_75t_R ALU___U240 ( .A(ALU__n1182), .B(ALU__n1184), .C(ALU__n1183), .Y(ALU__N371) );
  OA22x2_ASAP7_75t_R ALU___U245 ( .A1(ALU__n1336), .A2(ALU__n1485), .B1(ALU__n752), .B2(
        n925), .Y(ALU__n236) );
  OA221x2_ASAP7_75t_R ALU___U246 ( .A1(ALU__n1336), .A2(ALU__n1437), .B1(ALU__n1480), .B2(
        n925), .C(ALU__n1593), .Y(ALU__n235) );
  OR3x1_ASAP7_75t_R ALU___U247 ( .A(ALU__n1060), .B(ALU__n1062), .C(ALU__n1061), .Y(ALU__N370) );
  AO22x1_ASAP7_75t_R ALU___U250 ( .A1(ALU__N305), .A2(ALU__n1516), .B1(ALU__N337), .B2(ALU__n1504), .Y(
        n238) );
  OA22x2_ASAP7_75t_R ALU___U252 ( .A1(ALU__n1337), .A2(ALU__n1485), .B1(ALU__n751), .B2(
        n969), .Y(ALU__n242) );
  OA221x2_ASAP7_75t_R ALU___U253 ( .A1(ALU__n1337), .A2(ALU__n1438), .B1(ALU__n1473), .B2(
        n969), .C(ALU__n1591), .Y(ALU__n241) );
  OR3x1_ASAP7_75t_R ALU___U254 ( .A(ALU__n1117), .B(ALU__n1119), .C(ALU__n1118), .Y(ALU__N369) );
  AO22x1_ASAP7_75t_R ALU___U257 ( .A1(ALU__N304), .A2(ALU__n1516), .B1(ALU__N336), .B2(ALU__n1504), .Y(
        n244) );
  OA22x2_ASAP7_75t_R ALU___U259 ( .A1(ALU__n1014), .A2(ALU__n1486), .B1(ALU__n1123), .B2(
        n1020), .Y(ALU__n248) );
  OA221x2_ASAP7_75t_R ALU___U260 ( .A1(ALU__n1014), .A2(ALU__n1438), .B1(ALU__n1476), .B2(
        n1020), .C(ALU__n1600), .Y(ALU__n247) );
  OR3x1_ASAP7_75t_R ALU___U261 ( .A(ALU__n1094), .B(ALU__n1096), .C(ALU__n1095), .Y(ALU__N368) );
  AO22x1_ASAP7_75t_R ALU___U264 ( .A1(ALU__N303), .A2(ALU__n1516), .B1(ALU__N335), .B2(ALU__n1504), .Y(
        n250) );
  OA22x2_ASAP7_75t_R ALU___U266 ( .A1(ALU__n982), .A2(ALU__n1486), .B1(ALU__n1463), .B2(
        n1109), .Y(ALU__n254) );
  OA221x2_ASAP7_75t_R ALU___U267 ( .A1(ALU__n982), .A2(ALU__n1439), .B1(ALU__n1487), .B2(
        n1109), .C(ALU__n1592), .Y(ALU__n253) );
  OR3x1_ASAP7_75t_R ALU___U268 ( .A(ALU__n1138), .B(ALU__n1140), .C(ALU__n1139), .Y(ALU__N367) );
  OA22x2_ASAP7_75t_R ALU___U273 ( .A1(ALU__n1753), .A2(ALU__n1486), .B1(ALU__n1463), .B2(
        n1152), .Y(ALU__n260) );
  OA221x2_ASAP7_75t_R ALU___U274 ( .A1(ALU__n1753), .A2(ALU__n1439), .B1(ALU__n1471), .B2(
        n1152), .C(ALU__n1593), .Y(ALU__n259) );
  OR3x1_ASAP7_75t_R ALU___U275 ( .A(ALU__n1219), .B(ALU__n1221), .C(ALU__n1220), .Y(ALU__N366) );
  AO22x1_ASAP7_75t_R ALU___U278 ( .A1(ALU__N301), .A2(ALU__n1516), .B1(ALU__N333), .B2(ALU__n1504), .Y(
        n262) );
  OA22x2_ASAP7_75t_R ALU___U280 ( .A1(ALU__n1386), .A2(ALU__n1487), .B1(ALU__n1454), .B2(
        n1229), .Y(ALU__n266) );
  OA221x2_ASAP7_75t_R ALU___U281 ( .A1(ALU__n1386), .A2(ALU__ALU__n1445), .B1(ALU__n14), .B2(
        n1229), .C(ALU__n1592), .Y(ALU__n265) );
  OR3x1_ASAP7_75t_R ALU___U282 ( .A(ALU__n1146), .B(ALU__n1148), .C(ALU__n1147), .Y(ALU__N365) );
  AO22x1_ASAP7_75t_R ALU___U285 ( .A1(ALU__N300), .A2(ALU__n1515), .B1(ALU__N332), .B2(ALU__n1503), .Y(
        n268) );
  OA22x2_ASAP7_75t_R ALU___U287 ( .A1(ALU__n1389), .A2(ALU__n1487), .B1(ALU__n1460), .B2(
        n1029), .Y(ALU__n272) );
  OA221x2_ASAP7_75t_R ALU___U288 ( .A1(ALU__n1389), .A2(ALU__n1445), .B1(ALU__n1474), .B2(
        n1029), .C(ALU__n1589), .Y(ALU__n271) );
  OR3x1_ASAP7_75t_R ALU___U289 ( .A(ALU__n931), .B(ALU__n933), .C(ALU__n932), .Y(ALU__N364) );
  AO22x1_ASAP7_75t_R ALU___U292 ( .A1(ALU__N299), .A2(ALU__n1515), .B1(ALU__N331), .B2(ALU__n1503), .Y(
        n274) );
  OA22x2_ASAP7_75t_R ALU___U294 ( .A1(ALU__n1390), .A2(ALU__n1487), .B1(ALU__n1460), .B2(
        n929), .Y(ALU__n278) );
  OA221x2_ASAP7_75t_R ALU___U295 ( .A1(ALU__n1390), .A2(ALU__n1440), .B1(ALU__n1472), .B2(
        n929), .C(ALU__n1591), .Y(ALU__n277) );
  OR3x1_ASAP7_75t_R ALU___U296 ( .A(ALU__n1186), .B(ALU__n1188), .C(ALU__n1187), .Y(ALU__N363) );
  AO22x1_ASAP7_75t_R ALU___U299 ( .A1(ALU__N298), .A2(ALU__n1515), .B1(ALU__N330), .B2(ALU__n1503), .Y(
        n280) );
  OA22x2_ASAP7_75t_R ALU___U301 ( .A1(ALU__n1275), .A2(ALU__n1488), .B1(ALU__n1043), .B2(
        n1114), .Y(ALU__n284) );
  OA221x2_ASAP7_75t_R ALU___U302 ( .A1(ALU__n1275), .A2(ALU__n1440), .B1(ALU__n1474), .B2(
        n1114), .C(ALU__n1590), .Y(ALU__n283) );
  OR3x1_ASAP7_75t_R ALU___U303 ( .A(ALU__n962), .B(ALU__n964), .C(ALU__n963), .Y(ALU__N362) );
  AO22x1_ASAP7_75t_R ALU___U306 ( .A1(ALU__N297), .A2(ALU__n1515), .B1(ALU__N329), .B2(ALU__n1503), .Y(
        n286) );
  OA22x2_ASAP7_75t_R ALU___U308 ( .A1(ALU__n1363), .A2(ALU__n1488), .B1(ALU__n1042), .B2(
        n973), .Y(ALU__n290) );
  OA221x2_ASAP7_75t_R ALU___U309 ( .A1(ALU__n1363), .A2(ALU__n1441), .B1(ALU__n1473), .B2(
        n973), .C(ALU__n1592), .Y(ALU__n289) );
  OR3x1_ASAP7_75t_R ALU___U310 ( .A(ALU__n1268), .B(ALU__n1270), .C(ALU__n1269), .Y(ALU__N361) );
  AO22x1_ASAP7_75t_R ALU___U313 ( .A1(ALU__N296), .A2(ALU__n1515), .B1(ALU__N328), .B2(ALU__n1503), .Y(
        n292) );
  OA22x2_ASAP7_75t_R ALU___U315 ( .A1(ALU__n1387), .A2(ALU__n1488), .B1(ALU__n1041), .B2(
        n1233), .Y(ALU__n296) );
  OA221x2_ASAP7_75t_R ALU___U316 ( .A1(ALU__n1387), .A2(ALU__n1441), .B1(ALU__n1471), .B2(
        n1233), .C(ALU__n1587), .Y(ALU__n295) );
  OR3x1_ASAP7_75t_R ALU___U317 ( .A(ALU__n1223), .B(ALU__n1225), .C(ALU__n1224), .Y(ALU__N360) );
  AO22x1_ASAP7_75t_R ALU___U320 ( .A1(ALU__N295), .A2(ALU__n1515), .B1(ALU__N327), .B2(ALU__n1503), .Y(
        n298) );
  OA22x2_ASAP7_75t_R ALU___U322 ( .A1(ALU__n1360), .A2(ALU__n1489), .B1(ALU__n1104), .B2(
        n1174), .Y(ALU__n302) );
  OA221x2_ASAP7_75t_R ALU___U323 ( .A1(ALU__n1360), .A2(ALU__n1442), .B1(ALU__n1472), .B2(
        n1174), .C(ALU__n1593), .Y(ALU__n301) );
  OR3x1_ASAP7_75t_R ALU___U324 ( .A(ALU__n1142), .B(ALU__n1144), .C(ALU__n1143), .Y(ALU__N359) );
  AO22x1_ASAP7_75t_R ALU___U327 ( .A1(ALU__N294), .A2(ALU__n1514), .B1(ALU__N326), .B2(ALU__n1502), .Y(
        n304) );
  OA22x2_ASAP7_75t_R ALU___U329 ( .A1(ALU__n1421), .A2(ALU__n1489), .B1(ALU__n1103), .B2(
        n1060), .Y(ALU__n308) );
  OA221x2_ASAP7_75t_R ALU___U330 ( .A1(ALU__n1421), .A2(ALU__n1442), .B1(ALU__n1471), .B2(
        n1060), .C(ALU__n1587), .Y(ALU__n307) );
  OR3x1_ASAP7_75t_R ALU___U331 ( .A(ALU__n1000), .B(ALU__n1002), .C(ALU__n1001), .Y(ALU__N358) );
  AO22x1_ASAP7_75t_R ALU___U334 ( .A1(ALU__N293), .A2(ALU__n1514), .B1(ALU__N325), .B2(ALU__n1502), .Y(
        n310) );
  OA22x2_ASAP7_75t_R ALU___U336 ( .A1(ALU__n1301), .A2(ALU__n1489), .B1(ALU__n1102), .B2(ALU__n1032), 
        .Y(ALU__n314) );
  OA221x2_ASAP7_75t_R ALU___U337 ( .A1(ALU__n1301), .A2(ALU__n1443), .B1(ALU__n1469), .B2(ALU__n1032), 
        .C(ALU__n1588), .Y(ALU__n313) );
  OR3x1_ASAP7_75t_R ALU___U338 ( .A(ALU__n1098), .B(ALU__n1100), .C(ALU__n1099), .Y(ALU__N357) );
  AO22x1_ASAP7_75t_R ALU___U341 ( .A1(ALU__N292), .A2(ALU__n1514), .B1(ALU__N324), .B2(ALU__n1502), .Y(
        n316) );
  OA22x2_ASAP7_75t_R ALU___U343 ( .A1(ALU__n1415), .A2(ALU__n1490), .B1(ALU__n1463), .B2(
        n1015), .Y(ALU__n320) );
  OA221x2_ASAP7_75t_R ALU___U344 ( .A1(ALU__n1415), .A2(ALU__n1443), .B1(ALU__n1480), .B2(
        n1015), .C(ALU__n1587), .Y(ALU__n319) );
  OA221x2_ASAP7_75t_R ALU___U346 ( .A1(ALU__n1083), .A2(ALU__n1623), .B1(ALU__n1372), .B2(ALU__n1594), 
        .C(ALU__n1021), .Y(ALU__n323) );
  OA222x2_ASAP7_75t_R ALU___U348 ( .A1(ALU__n644), .A2(ALU__n1700), .B1(ALU__n1047), .B2(ALU__n1309), 
        .C1(n892), .C2(ALU__n582), .Y(ALU__n322) );
  OA22x2_ASAP7_75t_R ALU___U349 ( .A1(ALU__n1372), .A2(ALU__n1490), .B1(ALU__n1463), .B2(
        n964), .Y(ALU__n328) );
  MAJx2_ASAP7_75t_R ALU___U350 ( .A(n1091), .B(ALU__n1049), .C(ALU__n1308), .Y(ALU__n326) );
  OA221x2_ASAP7_75t_R ALU___U351 ( .A1(ALU__n1372), .A2(ALU__n1444), .B1(ALU__n1479), .B2(
        n964), .C(ALU__n1591), .Y(ALU__n325) );
  AND2x2_ASAP7_75t_R ALU___U355 ( .A(ALU__n668), .B(ALU_ctl[3]), .Y(ALU__n135) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW_rash_0___U3 ( .A(ALU_DW_rash_0__n687), .Y(ALU_DW_rash_0__n1) );
  INVxp33_ASAP7_75t_R ALU___ALU_DW_rash_0___U4 ( .A(ALU_DW_rash_0__n2), .Y(ALU_DW_rash_0__n687) );
  NOR2x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U5 ( .A(ALU_DW_rash_0__n285), .B(ALU_DW_rash_0__n4), .Y(ALU_DW_rash_0__n3) );
  NOR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U6 ( .A(ALU_DW_rash_0__n456), .B(ALU_DW_rash_0__n183), .Y(ALU_DW_rash_0__n5) );
  NOR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U7 ( .A(ALU_DW_rash_0__n428), .B(ALU_DW_rash_0__n395), .Y(ALU_DW_rash_0__n6) );
  NOR2xp67_ASAP7_75t_R ALU___ALU_DW_rash_0___U8 ( .A(ALU_DW_rash_0__n6), .B(ALU_DW_rash_0__n7), .Y(ALU_DW_rash_0__n2) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW_rash_0___U9 ( .A(ALU_DW_rash_0__n205), .B(ALU_DW_rash_0__n360), .Y(ALU_DW_rash_0__n8) );
  INVx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U10 ( .A(ALU_DW_rash_0__n8), .Y(ALU_DW_rash_0__n4) );
  NOR2x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U11 ( .A(ALU_DW_rash_0__n3), .B(ALU_DW_rash_0__n5), .Y(ALU_DW_rash_0__n9) );
  INVx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U12 ( .A(ALU_DW_rash_0__n9), .Y(ALU_DW_rash_0__n7) );
  CKINVDCx6p67_ASAP7_75t_R ALU___ALU_DW_rash_0___U13 ( .A(ALU_DW_rash_0__n236), .Y(ALU_DW_rash_0__n428) );
  CKINVDCx6p67_ASAP7_75t_R ALU___ALU_DW_rash_0___U14 ( .A(ALU_DW_rash_0__n228), .Y(ALU_DW_rash_0__n456) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U15 ( .A(ALU_DW_rash_0__n707), .Y(ALU_DW_rash_0__n10) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U16 ( .A(ALU_DW_rash_0__n178), .Y(ALU_DW_rash_0__n573) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U17 ( .A(ALU_DW_rash_0__n426), .Y(ALU_DW_rash_0__n28) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U18 ( .A(ALU_DW_rash_0__n706), .Y(ALU_DW_rash_0__n11) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U19 ( .A(ALU_DW_rash_0__n179), .Y(ALU_DW_rash_0__n572) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U20 ( .A(ALU_DW_rash_0__n709), .Y(ALU_DW_rash_0__n12) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U21 ( .A(ALU_DW_rash_0__n28), .Y(ALU_DW_rash_0__n379) );
  CKINVDCx6p67_ASAP7_75t_R ALU___ALU_DW_rash_0___U22 ( .A(ALU_DW_rash_0__n184), .Y(ALU_DW_rash_0__n497) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U23 ( .A(ALU_DW_rash_0__n22), .Y(ALU_DW_rash_0__n575) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U24 ( .A(ALU__n73), .Y(ALU_DW_rash_0__n13) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW_rash_0___U25 ( .A(ALU_DW_rash_0__n571), .Y(ALU_DW_rash_0__n14) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U26 ( .A(ALU_DW_rash_0__n571), .Y(ALU_DW_rash_0__n15) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW_rash_0___U27 ( .A(ALU_DW_rash_0__n25), .Y(ALU_DW_rash_0__n16) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U28 ( .A(ALU_DW_rash_0__n305), .Y(ALU_DW_rash_0__n25) );
  CKINVDCx20_ASAP7_75t_R ALU___ALU_DW_rash_0___U29 ( .A(ALU_DW_rash_0__n19), .Y(ALU_DW_rash_0__n17) );
  CKINVDCx20_ASAP7_75t_R ALU___ALU_DW_rash_0___U30 ( .A(ALU_DW_rash_0__n17), .Y(ALU_DW_rash_0__n18) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW_rash_0___U31 ( .A(ALU_DW_rash_0__n201), .Y(ALU_DW_rash_0__n19) );
  CKINVDCx20_ASAP7_75t_R ALU___ALU_DW_rash_0___U32 ( .A(ALU_DW_rash_0__n18), .Y(ALU_DW_rash_0__n517) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U33 ( .A(ALU_DW_rash_0__n202), .Y(ALU_DW_rash_0__n201) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U34 ( .A(ALU__n80), .Y(ALU_DW_rash_0__n20) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U35 ( .A(ALU__n348), .Y(ALU_DW_rash_0__n47) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U36 ( .A(ALU_DW_rash_0__n23), .Y(ALU_DW_rash_0__n21) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U37 ( .A(ALU_DW_rash_0__n24), .Y(ALU_DW_rash_0__n22) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U38 ( .A(ALU_DW_rash_0__n576), .Y(ALU_DW_rash_0__n23) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U39 ( .A(ALU_DW_rash_0__n23), .Y(ALU_DW_rash_0__n24) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U40 ( .A(ALU_DW_rash_0__n306), .Y(ALU_DW_rash_0__n305) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U41 ( .A(n1029), .Y(ALU_DW_rash_0__n26) );
  INVx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U42 ( .A(ALU_DW_rash_0__n57), .Y(ALU_DW_rash_0__n27) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U43 ( .A(ALU_DW_rash_0__n426), .Y(ALU_DW_rash_0__n29) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U44 ( .A(ALU_DW_rash_0__n426), .Y(ALU_DW_rash_0__n30) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U45 ( .A(ALU_DW_rash_0__n47), .Y(ALU_DW_rash_0__n308) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U46 ( .A(ALU_DW_rash_0__n561), .Y(ALU_DW_rash_0__n297) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U47 ( .A(ALU_DW_rash_0__n33), .Y(ALU_DW_rash_0__n31) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U48 ( .A(ALU_DW_rash_0__n33), .Y(ALU_DW_rash_0__n32) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U49 ( .A(ALU_DW_rash_0__n39), .Y(ALU_DW_rash_0__n33) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U50 ( .A(ALU_DW_rash_0__n37), .Y(ALU_DW_rash_0__n34) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U51 ( .A(ALU_DW_rash_0__n341), .Y(ALU_DW_rash_0__n35) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U52 ( .A(ALU_DW_rash_0__n28), .Y(ALU_DW_rash_0__n380) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U53 ( .A(ALU_DW_rash_0__n56), .Y(ALU_DW_rash_0__n36) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U54 ( .A(ALU_DW_rash_0__n308), .Y(ALU_DW_rash_0__n599) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U55 ( .A(ALU_DW_rash_0__n624), .Y(ALU_DW_rash_0__n37) );
  CKINVDCx10_ASAP7_75t_R ALU___ALU_DW_rash_0___U56 ( .A(ALU_DW_rash_0__n283), .Y(ALU_DW_rash_0__n454) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U57 ( .A(ALU_DW_rash_0__n241), .Y(ALU_DW_rash_0__n240) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U58 ( .A(ALU_DW_rash_0__n34), .Y(ALU_DW_rash_0__n241) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U59 ( .A(n1020), .Y(ALU_DW_rash_0__n38) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U60 ( .A(ALU_DW_rash_0__n574), .Y(ALU_DW_rash_0__n39) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U61 ( .A(ALU_DW_rash_0__n45), .Y(ALU_DW_rash_0__n40) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U62 ( .A(ALU_DW_rash_0__n642), .Y(ALU_DW_rash_0__n41) );
  CKINVDCx9p33_ASAP7_75t_R ALU___ALU_DW_rash_0___U63 ( .A(ALU_DW_rash_0__n108), .Y(ALU_DW_rash_0__n410) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U64 ( .A(ALU_DW_rash_0__n43), .Y(ALU_DW_rash_0__n42) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U65 ( .A(ALU_DW_rash_0__n612), .Y(ALU_DW_rash_0__n43) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U66 ( .A(ALU_DW_rash_0__n116), .Y(ALU_DW_rash_0__n44) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U67 ( .A(ALU_DW_rash_0__n630), .Y(ALU_DW_rash_0__n45) );
  CKINVDCx10_ASAP7_75t_R ALU___ALU_DW_rash_0___U68 ( .A(ALU_DW_rash_0__n414), .Y(ALU_DW_rash_0__n466) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U69 ( .A(ALU_DW_rash_0__n436), .Y(ALU_DW_rash_0__n435) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U70 ( .A(ALU_DW_rash_0__n40), .Y(ALU_DW_rash_0__n436) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U71 ( .A(ALU_DW_rash_0__n62), .Y(ALU_DW_rash_0__n46) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U72 ( .A(ALU__n348), .Y(ALU_DW_rash_0__n48) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U73 ( .A(ALU__n348), .Y(ALU_DW_rash_0__n49) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U74 ( .A(ALU_DW_rash_0__n583), .Y(ALU_DW_rash_0__n50) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U75 ( .A(ALU_DW_rash_0__n583), .Y(ALU_DW_rash_0__n51) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U76 ( .A(ALU_DW_rash_0__n66), .Y(ALU_DW_rash_0__n52) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U77 ( .A(ALU_DW_rash_0__n66), .Y(ALU_DW_rash_0__n53) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U78 ( .A(ALU_DW_rash_0__n36), .Y(ALU_DW_rash_0__n54) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U79 ( .A(ALU_DW_rash_0__n36), .Y(ALU_DW_rash_0__n55) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U80 ( .A(ALU_DW_rash_0__n304), .Y(ALU_DW_rash_0__n56) );
  INVx5_ASAP7_75t_R ALU___ALU_DW_rash_0___U81 ( .A(ALU_DW_rash_0__n54), .Y(ALU_DW_rash_0__n563) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U82 ( .A(ALU_DW_rash_0__n178), .Y(ALU_DW_rash_0__n304) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U83 ( .A(ALU_DW_rash_0__n306), .Y(ALU_DW_rash_0__n307) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U84 ( .A(ALU_DW_rash_0__n662), .Y(ALU_DW_rash_0__n57) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U85 ( .A(ALU_DW_rash_0__n539), .Y(ALU_DW_rash_0__n58) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U86 ( .A(ALU_DW_rash_0__n539), .Y(ALU_DW_rash_0__n59) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U87 ( .A(ALU_DW_rash_0__n539), .Y(ALU_DW_rash_0__n60) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U88 ( .A(ALU_DW_rash_0__n58), .B(ALU_DW_rash_0__n380), .Y(ALU_DW_rash_0__n601) );
  CKINVDCx14_ASAP7_75t_R ALU___ALU_DW_rash_0___U89 ( .A(ALU_DW_rash_0__n343), .Y(ALU_DW_rash_0__n539) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U90 ( .A(ALU_DW_rash_0__n653), .Y(ALU_DW_rash_0__n61) );
  CKINVDCx11_ASAP7_75t_R ALU___ALU_DW_rash_0___U91 ( .A(ALU_DW_rash_0__n511), .Y(ALU_DW_rash_0__n585) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U92 ( .A(ALU_DW_rash_0__n176), .Y(ALU_DW_rash_0__n584) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U93 ( .A(ALU_DW_rash_0__n73), .Y(ALU_DW_rash_0__n403) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U94 ( .A(ALU_DW_rash_0__n633), .Y(ALU_DW_rash_0__n62) );
  CKINVDCx10_ASAP7_75t_R ALU___ALU_DW_rash_0___U95 ( .A(ALU_DW_rash_0__n238), .Y(ALU_DW_rash_0__n477) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U96 ( .A(ALU_DW_rash_0__n327), .Y(ALU_DW_rash_0__n326) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U97 ( .A(ALU_DW_rash_0__n46), .Y(ALU_DW_rash_0__n327) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U98 ( .A(ALU_DW_rash_0__n130), .Y(ALU_DW_rash_0__n63) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U99 ( .A(ALU_DW_rash_0__n623), .Y(ALU_DW_rash_0__n64) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U100 ( .A1(ALU_DW_rash_0__n554), .A2(ALU_DW_rash_0__n434), .B1(ALU_DW_rash_0__n564), .B2(n973), .C(
        n374), .Y(ALU_DW_rash_0__n623) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U101 ( .A(ALU_DW_rash_0__n735), .Y(ALU_DW_rash_0__n65) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U102 ( .A(ALU_DW_rash_0__n529), .Y(ALU_DW_rash_0__n526) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U103 ( .A(ALU_DW_rash_0__n50), .Y(ALU_DW_rash_0__n580) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U104 ( .A(ALU_DW_rash_0__n101), .Y(ALU_DW_rash_0__n66) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U105 ( .A(ALU__n368), .Y(ALU_DW_rash_0__n67) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U106 ( .A(ALU_DW_rash_0__n639), .Y(ALU_DW_rash_0__n68) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U107 ( .A(ALU_DW_rash_0__n115), .Y(ALU_DW_rash_0__n69) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U108 ( .A(ALU_DW_rash_0__n629), .Y(ALU_DW_rash_0__n70) );
  INVx5_ASAP7_75t_R ALU___ALU_DW_rash_0___U109 ( .A(ALU_DW_rash_0__n481), .Y(ALU_DW_rash_0__n550) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U110 ( .A1(ALU_DW_rash_0__n550), .A2(n973), .B1(ALU_DW_rash_0__n570), .B2(n1233), .C(
        n416), .Y(ALU_DW_rash_0__n629) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U111 ( .A(ALU_DW_rash_0__n739), .Y(ALU_DW_rash_0__n71) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U112 ( .A(ALU_DW_rash_0__n97), .Y(ALU_DW_rash_0__n590) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U113 ( .A(ALU_DW_rash_0__n96), .Y(ALU_DW_rash_0__n589) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U114 ( .A(ALU_DW_rash_0__n646), .Y(ALU_DW_rash_0__n72) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW_rash_0___U115 ( .A(ALU_DW_rash_0__n140), .Y(ALU_DW_rash_0__n73) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U116 ( .A(ALU_DW_rash_0__n141), .Y(ALU_DW_rash_0__n74) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U117 ( .A(ALU_DW_rash_0__n74), .Y(ALU_DW_rash_0__n140) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U118 ( .A(ALU_DW_rash_0__n671), .Y(ALU_DW_rash_0__n75) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U119 ( .A(ALU_DW_rash_0__n314), .Y(ALU_DW_rash_0__n452) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U120 ( .A(ALU_DW_rash_0__n737), .Y(ALU_DW_rash_0__n76) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U121 ( .A(ALU_DW_rash_0__n743), .Y(ALU_DW_rash_0__n77) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U122 ( .A(ALU_DW_rash_0__n79), .Y(ALU_DW_rash_0__n78) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U123 ( .A(ALU_DW_rash_0__n621), .Y(ALU_DW_rash_0__n79) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U124 ( .A(ALU_DW_rash_0__n94), .Y(ALU_DW_rash_0__n80) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U125 ( .A1(ALU_DW_rash_0__n552), .A2(n1109), .B1(ALU_DW_rash_0__n566), .B2(ALU_DW_rash_0__n470), .C(
        n394), .Y(ALU_DW_rash_0__n621) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U126 ( .A(ALU_DW_rash_0__n82), .Y(ALU_DW_rash_0__n81) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U127 ( .A(ALU_DW_rash_0__n703), .Y(ALU_DW_rash_0__n82) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U128 ( .A(ALU_DW_rash_0__n84), .Y(ALU_DW_rash_0__n83) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U129 ( .A(ALU_DW_rash_0__n602), .Y(ALU_DW_rash_0__n84) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U130 ( .A(ALU_DW_rash_0__n383), .Y(ALU_DW_rash_0__n85) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U131 ( .A(ALU_DW_rash_0__n383), .Y(ALU_DW_rash_0__n86) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U132 ( .A(ALU_DW_rash_0__n169), .Y(ALU_DW_rash_0__n87) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U133 ( .A(ALU_DW_rash_0__n632), .Y(ALU_DW_rash_0__n88) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U134 ( .A1(ALU_DW_rash_0__n554), .A2(n1233), .B1(ALU_DW_rash_0__n568), .B2(ALU_DW_rash_0__n342), .C(
        n391), .Y(ALU_DW_rash_0__n632) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U135 ( .A(ALU_DW_rash_0__n741), .Y(ALU_DW_rash_0__n89) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U136 ( .A(ALU_DW_rash_0__n652), .Y(ALU_DW_rash_0__n90) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U137 ( .A(ALU_DW_rash_0__n92), .Y(ALU_DW_rash_0__n91) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U138 ( .A(ALU_DW_rash_0__n627), .Y(ALU_DW_rash_0__n92) );
  INVx5_ASAP7_75t_R ALU___ALU_DW_rash_0___U139 ( .A(ALU_DW_rash_0__n522), .Y(ALU_DW_rash_0__n554) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U140 ( .A1(ALU_DW_rash_0__n554), .A2(ALU_DW_rash_0__n471), .B1(ALU_DW_rash_0__n567), .B2(ALU_DW_rash_0__n199), .C(
        n422), .Y(ALU_DW_rash_0__n627) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U141 ( .A(ALU__n410), .Y(ALU_DW_rash_0__n93) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U142 ( .A(ALU_DW_rash_0__n95), .Y(ALU_DW_rash_0__n94) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U143 ( .A(ALU_DW_rash_0__n78), .Y(ALU_DW_rash_0__n95) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U144 ( .A(ALU_DW_rash_0__n80), .Y(ALU_DW_rash_0__n393) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U145 ( .A(ALU_DW_rash_0__n98), .Y(ALU_DW_rash_0__n96) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U146 ( .A(ALU_DW_rash_0__n98), .Y(ALU_DW_rash_0__n97) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U147 ( .A(ALU_DW_rash_0__n535), .Y(ALU_DW_rash_0__n98) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U148 ( .A(ALU_DW_rash_0__n53), .Y(ALU_DW_rash_0__n99) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U149 ( .A(ALU_DW_rash_0__n52), .Y(ALU_DW_rash_0__n100) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U150 ( .A(ALU_DW_rash_0__n558), .Y(ALU_DW_rash_0__n101) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U151 ( .A(ALU_DW_rash_0__n47), .Y(ALU_DW_rash_0__n310) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U152 ( .A(ALU_DW_rash_0__n103), .Y(ALU_DW_rash_0__n102) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U153 ( .A(ALU_DW_rash_0__n514), .Y(ALU_DW_rash_0__n103) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U154 ( .A(ALU_DW_rash_0__n102), .Y(ALU_DW_rash_0__n104) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U155 ( .A(ALU_DW_rash_0__n102), .Y(ALU_DW_rash_0__n200) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U156 ( .A(ALU_DW_rash_0__n490), .Y(ALU_DW_rash_0__n105) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U157 ( .A(ALU_DW_rash_0__n490), .Y(ALU_DW_rash_0__n106) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U158 ( .A(ALU_DW_rash_0__n742), .Y(ALU_DW_rash_0__n107) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW_rash_0___U159 ( .A(ALU_DW_rash_0__n109), .Y(ALU_DW_rash_0__n108) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U160 ( .A(ALU_DW_rash_0__n41), .Y(ALU_DW_rash_0__n109) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U161 ( .A(ALU_DW_rash_0__n740), .Y(ALU_DW_rash_0__n110) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U162 ( .A(ALU_DW_rash_0__n677), .Y(ALU_DW_rash_0__n111) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U163 ( .A(ALU_DW_rash_0__n113), .Y(ALU_DW_rash_0__n112) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U164 ( .A(ALU_DW_rash_0__n664), .Y(ALU_DW_rash_0__n113) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U165 ( .A1(ALU_DW_rash_0__n551), .A2(n920), .B1(ALU_DW_rash_0__n565), .B2(n1160), .C(
        n404), .Y(ALU_DW_rash_0__n664) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U166 ( .A(ALU_DW_rash_0__n69), .Y(ALU_DW_rash_0__n114) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U167 ( .A(ALU_DW_rash_0__n70), .Y(ALU_DW_rash_0__n115) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U168 ( .A(ALU_DW_rash_0__n114), .Y(ALU_DW_rash_0__n418) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U169 ( .A(ALU_DW_rash_0__n117), .Y(ALU_DW_rash_0__n116) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U170 ( .A(ALU_DW_rash_0__n91), .Y(ALU_DW_rash_0__n117) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U171 ( .A(ALU_DW_rash_0__n44), .Y(ALU_DW_rash_0__n424) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U172 ( .A(ALU_DW_rash_0__n119), .Y(ALU_DW_rash_0__n118) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U173 ( .A(ALU_DW_rash_0__n635), .Y(ALU_DW_rash_0__n119) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U174 ( .A1(ALU_DW_rash_0__n342), .A2(ALU_DW_rash_0__n552), .B1(n1060), .B2(ALU_DW_rash_0__n564), .C(
        n431), .Y(ALU_DW_rash_0__n635) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U175 ( .A(ALU_DW_rash_0__n736), .Y(ALU_DW_rash_0__n120) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U176 ( .A(ALU_DW_rash_0__n122), .Y(ALU_DW_rash_0__n121) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U177 ( .A(ALU_DW_rash_0__n618), .Y(ALU_DW_rash_0__n122) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U178 ( .A(ALU_DW_rash_0__n124), .Y(ALU_DW_rash_0__n123) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U179 ( .A(ALU_DW_rash_0__n651), .Y(ALU_DW_rash_0__n124) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U180 ( .A(ALU_DW_rash_0__n126), .Y(ALU_DW_rash_0__n125) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U181 ( .A(ALU_DW_rash_0__n650), .Y(ALU_DW_rash_0__n126) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U182 ( .A1(n1060), .A2(ALU_DW_rash_0__n551), .B1(ALU_DW_rash_0__n405), .B2(ALU_DW_rash_0__n570), .C(
        n242), .Y(ALU_DW_rash_0__n650) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U183 ( .A(ALU_DW_rash_0__n710), .Y(ALU_DW_rash_0__n127) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U184 ( .A(ALU_DW_rash_0__n744), .Y(ALU_DW_rash_0__n128) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U185 ( .A(ALU_DW_rash_0__n398), .B(ALU_DW_rash_0__n58), .Y(ALU_DW_rash_0__n679) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U186 ( .A(ALU_DW_rash_0__n63), .Y(ALU_DW_rash_0__n129) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U187 ( .A(ALU_DW_rash_0__n64), .Y(ALU_DW_rash_0__n130) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U188 ( .A(ALU_DW_rash_0__n129), .Y(ALU_DW_rash_0__n376) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U189 ( .A(ALU_DW_rash_0__n132), .Y(ALU_DW_rash_0__n131) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U190 ( .A(ALU_DW_rash_0__n669), .Y(ALU_DW_rash_0__n132) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U191 ( .A(ALU_DW_rash_0__n134), .Y(ALU_DW_rash_0__n133) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U192 ( .A(ALU_DW_rash_0__n668), .Y(ALU_DW_rash_0__n134) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U193 ( .A1(ALU_DW_rash_0__n406), .A2(ALU_DW_rash_0__n555), .B1(n1015), .B2(ALU_DW_rash_0__n567), .C(
        n229), .Y(ALU_DW_rash_0__n668) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW_rash_0___U194 ( .A(ALU_DW_rash_0__n235), .Y(ALU_DW_rash_0__n225) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U195 ( .A(ALU_DW_rash_0__n745), .Y(ALU_DW_rash_0__n135) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U196 ( .A(ALU_DW_rash_0__n137), .Y(ALU_DW_rash_0__n136) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U197 ( .A(ALU_DW_rash_0__n617), .Y(ALU_DW_rash_0__n137) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U198 ( .A1(ALU_DW_rash_0__n553), .A2(n929), .B1(ALU_DW_rash_0__n563), .B2(ALU_DW_rash_0__n434), .C(
        n361), .Y(ALU_DW_rash_0__n617) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U199 ( .A(ALU_DW_rash_0__n139), .Y(ALU_DW_rash_0__n138) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U200 ( .A(ALU_DW_rash_0__n90), .Y(ALU_DW_rash_0__n139) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U201 ( .A(ALU_DW_rash_0__n170), .Y(ALU_DW_rash_0__n507) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U202 ( .A(ALU_DW_rash_0__n112), .Y(ALU_DW_rash_0__n141) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U203 ( .A(ALU_DW_rash_0__n143), .Y(ALU_DW_rash_0__n142) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U204 ( .A(ALU_DW_rash_0__n700), .Y(ALU_DW_rash_0__n143) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U205 ( .A(ALU_DW_rash_0__n145), .Y(ALU_DW_rash_0__n144) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U206 ( .A(ALU_DW_rash_0__n701), .Y(ALU_DW_rash_0__n145) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U207 ( .A1(n1015), .A2(ALU_DW_rash_0__n554), .B1(n964), .B2(ALU_DW_rash_0__n568), .C(
        n211), .Y(ALU_DW_rash_0__n700) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW_rash_0___U208 ( .A(ALU_DW_rash_0__n180), .Y(ALU_DW_rash_0__n146) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U209 ( .A(ALU_DW_rash_0__n181), .Y(ALU_DW_rash_0__n180) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U210 ( .A(ALU_DW_rash_0__n515), .Y(ALU_DW_rash_0__n147) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U211 ( .A(ALU_DW_rash_0__n515), .Y(ALU_DW_rash_0__n148) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U212 ( .A(ALU_DW_rash_0__n515), .Y(ALU_DW_rash_0__n149) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U213 ( .A(n1073), .Y(ALU_DW_rash_0__n150) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U214 ( .A(ALU_DW_rash_0__n670), .Y(ALU_DW_rash_0__n151) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U215 ( .A(ALU_DW_rash_0__n153), .Y(ALU_DW_rash_0__n152) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U216 ( .A(ALU_DW_rash_0__n136), .Y(ALU_DW_rash_0__n153) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U217 ( .A(ALU_DW_rash_0__n155), .Y(ALU_DW_rash_0__n154) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U218 ( .A(ALU_DW_rash_0__n42), .Y(ALU_DW_rash_0__n155) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U219 ( .A(ALU_DW_rash_0__n157), .Y(ALU_DW_rash_0__n156) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U220 ( .A(ALU_DW_rash_0__n665), .Y(ALU_DW_rash_0__n157) );
  CKINVDCx5p33_ASAP7_75t_R ALU___ALU_DW_rash_0___U221 ( .A(ALU_DW_rash_0__n156), .Y(ALU_DW_rash_0__n440) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U222 ( .A(ALU_DW_rash_0__n159), .Y(ALU_DW_rash_0__n158) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U223 ( .A(ALU_DW_rash_0__n659), .Y(ALU_DW_rash_0__n159) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U224 ( .A(ALU_DW_rash_0__n338), .Y(ALU_DW_rash_0__n160) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U225 ( .A(ALU_DW_rash_0__n162), .Y(ALU_DW_rash_0__n161) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U226 ( .A(ALU_DW_rash_0__n643), .Y(ALU_DW_rash_0__n162) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U227 ( .A(ALU_DW_rash_0__n165), .Y(ALU_DW_rash_0__n163) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U228 ( .A(ALU_DW_rash_0__n166), .Y(ALU_DW_rash_0__n164) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U229 ( .A(ALU_DW_rash_0__n106), .Y(ALU_DW_rash_0__n165) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U230 ( .A(ALU_DW_rash_0__n105), .Y(ALU_DW_rash_0__n166) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U231 ( .A(ALU_DW_rash_0__n360), .B(ALU_DW_rash_0__n597), .Y(ALU_DW_rash_0__n643) );
  CKINVDCx9p33_ASAP7_75t_R ALU___ALU_DW_rash_0___U232 ( .A(ALU_DW_rash_0__n225), .Y(ALU_DW_rash_0__n597) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U233 ( .A(ALU_DW_rash_0__n161), .Y(ALU_DW_rash_0__n490) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U234 ( .A(ALU_DW_rash_0__n398), .Y(ALU_DW_rash_0__n167) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U235 ( .A(ALU_DW_rash_0__n87), .Y(ALU_DW_rash_0__n168) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U236 ( .A(ALU_DW_rash_0__n88), .Y(ALU_DW_rash_0__n169) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U237 ( .A(ALU_DW_rash_0__n168), .Y(ALU_DW_rash_0__n390) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U238 ( .A(ALU_DW_rash_0__n171), .Y(ALU_DW_rash_0__n170) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U239 ( .A(ALU_DW_rash_0__n667), .Y(ALU_DW_rash_0__n171) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U240 ( .A(ALU_DW_rash_0__n636), .Y(ALU_DW_rash_0__n172) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U241 ( .A(ALU_DW_rash_0__n193), .Y(ALU_DW_rash_0__n173) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U242 ( .A(ALU_DW_rash_0__n193), .Y(ALU_DW_rash_0__n174) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U243 ( .A(ALU_DW_rash_0__n525), .Y(ALU_DW_rash_0__n175) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U244 ( .A(ALU_DW_rash_0__n177), .Y(ALU_DW_rash_0__n176) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U245 ( .A(ALU_DW_rash_0__n72), .Y(ALU_DW_rash_0__n177) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U246 ( .A(ALU_DW_rash_0__n32), .Y(ALU_DW_rash_0__n178) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U247 ( .A(ALU_DW_rash_0__n31), .Y(ALU_DW_rash_0__n179) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U248 ( .A(ALU_DW_rash_0__n21), .Y(ALU_DW_rash_0__n574) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U249 ( .A(ALU_DW_rash_0__n610), .Y(ALU_DW_rash_0__n181) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U250 ( .A(ALU_DW_rash_0__n531), .Y(ALU_DW_rash_0__n182) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U251 ( .A(ALU_DW_rash_0__n531), .Y(ALU_DW_rash_0__n183) );
  CKINVDCx9p33_ASAP7_75t_R ALU___ALU_DW_rash_0___U252 ( .A(ALU_DW_rash_0__n146), .Y(ALU_DW_rash_0__n531) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U253 ( .A(ALU_DW_rash_0__n185), .Y(ALU_DW_rash_0__n184) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U254 ( .A(ALU_DW_rash_0__n638), .Y(ALU_DW_rash_0__n185) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U255 ( .A(ALU_DW_rash_0__n187), .Y(ALU_DW_rash_0__n186) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U256 ( .A(ALU_DW_rash_0__n702), .Y(ALU_DW_rash_0__n187) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U257 ( .A(ALU_DW_rash_0__n498), .Y(ALU_DW_rash_0__n188) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U258 ( .A(ALU_DW_rash_0__n190), .Y(ALU_DW_rash_0__n189) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U259 ( .A(ALU_DW_rash_0__n704), .Y(ALU_DW_rash_0__n190) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U260 ( .A(ALU_DW_rash_0__n192), .Y(ALU_DW_rash_0__n191) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U261 ( .A(ALU_DW_rash_0__n705), .Y(ALU_DW_rash_0__n192) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U262 ( .A(ALU_DW_rash_0__n497), .B(ALU_DW_rash_0__n310), .Y(ALU_DW_rash_0__n658) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U263 ( .A(ALU_DW_rash_0__n592), .Y(ALU_DW_rash_0__n193) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U264 ( .A(ALU_DW_rash_0__n196), .Y(ALU_DW_rash_0__n194) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U265 ( .A(ALU_DW_rash_0__n196), .Y(ALU_DW_rash_0__n195) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U266 ( .A(ALU_DW_rash_0__n294), .Y(ALU_DW_rash_0__n196) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U267 ( .A(ALU_DW_rash_0__n556), .Y(ALU_DW_rash_0__n197) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U268 ( .A(ALU_DW_rash_0__n734), .Y(ALU_DW_rash_0__n198) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U269 ( .A(n1229), .Y(ALU_DW_rash_0__n199) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U270 ( .A(ALU_DW_rash_0__n55), .Y(ALU_DW_rash_0__n564) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U271 ( .A(ALU_DW_rash_0__n641), .Y(ALU_DW_rash_0__n202) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U272 ( .A(ALU_DW_rash_0__n603), .Y(ALU_DW_rash_0__n203) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U273 ( .A(ALU_DW_rash_0__n205), .Y(ALU_DW_rash_0__n204) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U274 ( .A(ALU_DW_rash_0__n167), .Y(ALU_DW_rash_0__n205) );
  OR2x4_ASAP7_75t_R ALU___ALU_DW_rash_0___U275 ( .A(ALU_DW_rash_0__n476), .B(ALU_DW_rash_0__n497), .Y(ALU_DW_rash_0__n603) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U276 ( .A(ALU_DW_rash_0__n207), .Y(ALU_DW_rash_0__n206) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U277 ( .A(ALU_DW_rash_0__n606), .Y(ALU_DW_rash_0__n207) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U278 ( .A(ALU_DW_rash_0__n209), .Y(ALU_DW_rash_0__n208) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U279 ( .A(ALU_DW_rash_0__n151), .Y(ALU_DW_rash_0__n209) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U280 ( .A(ALU_DW_rash_0__n281), .Y(ALU_DW_rash_0__n505) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U281 ( .A(ALU_DW_rash_0__n368), .Y(ALU_DW_rash_0__n495) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U282 ( .A(ALU_DW_rash_0__n666), .Y(ALU_DW_rash_0__n210) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U283 ( .A(ALU_DW_rash_0__n719), .Y(ALU_DW_rash_0__n211) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U284 ( .A(ALU_DW_rash_0__n142), .Y(ALU_DW_rash_0__n212) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U285 ( .A1(ALU_DW_rash_0__n309), .A2(ALU_DW_rash_0__n400), .B1(ALU_DW_rash_0__n320), .B2(ALU_DW_rash_0__n476), .Y(
        n701) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U286 ( .A(ALU_DW_rash_0__n144), .Y(ALU_DW_rash_0__n213) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U287 ( .A(ALU_DW_rash_0__n648), .Y(ALU_DW_rash_0__n214) );
  INVx5_ASAP7_75t_R ALU___ALU_DW_rash_0___U288 ( .A(ALU_DW_rash_0__n214), .Y(ALU_DW_rash_0__n492) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U289 ( .A(ALU_DW_rash_0__n216), .Y(ALU_DW_rash_0__n215) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U290 ( .A(ALU_DW_rash_0__n628), .Y(ALU_DW_rash_0__n216) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U291 ( .A(ALU_DW_rash_0__n215), .Y(ALU_DW_rash_0__n462) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U292 ( .A(ALU_DW_rash_0__n218), .Y(ALU_DW_rash_0__n217) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U293 ( .A(ALU_DW_rash_0__n614), .Y(ALU_DW_rash_0__n218) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U294 ( .A(ALU_DW_rash_0__n217), .Y(ALU_DW_rash_0__n464) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U295 ( .A(ALU_DW_rash_0__n637), .Y(ALU_DW_rash_0__n219) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U296 ( .A(ALU_DW_rash_0__n640), .Y(ALU_DW_rash_0__n220) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U297 ( .A(ALU_DW_rash_0__n118), .Y(ALU_DW_rash_0__n221) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U298 ( .A(ALU_DW_rash_0__n521), .Y(ALU_DW_rash_0__n552) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U299 ( .A1(ALU_DW_rash_0__n452), .A2(ALU_DW_rash_0__n458), .B1(ALU_DW_rash_0__n85), .B2(ALU_DW_rash_0__n204), .C(
        n223), .Y(ALU_DW_rash_0__n740) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U300 ( .A(ALU_DW_rash_0__n110), .Y(ALU__N300) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U301 ( .A(ALU_DW_rash_0__n224), .Y(ALU_DW_rash_0__n223) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U302 ( .A(ALU_DW_rash_0__n604), .Y(ALU_DW_rash_0__n224) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U303 ( .A(ALU_DW_rash_0__n227), .Y(ALU_DW_rash_0__n226) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U304 ( .A(ALU_DW_rash_0__n111), .Y(ALU_DW_rash_0__n227) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U305 ( .A(ALU_DW_rash_0__n620), .Y(ALU_DW_rash_0__n228) );
  CKINVDCx5p33_ASAP7_75t_R ALU___ALU_DW_rash_0___U306 ( .A(ALU_DW_rash_0__n355), .Y(ALU_DW_rash_0__n542) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U307 ( .A(ALU_DW_rash_0__n674), .Y(ALU_DW_rash_0__n229) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U308 ( .A1(ALU_DW_rash_0__n311), .A2(ALU_DW_rash_0__n449), .B1(ALU_DW_rash_0__n287), .B2(ALU_DW_rash_0__n476), .Y(
        n669) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U309 ( .A(ALU_DW_rash_0__n131), .Y(ALU_DW_rash_0__n230) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U310 ( .A(ALU_DW_rash_0__n133), .Y(ALU_DW_rash_0__n231) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U311 ( .A1(ALU_DW_rash_0__n376), .A2(ALU_DW_rash_0__n458), .B1(ALU_DW_rash_0__n240), .B2(ALU_DW_rash_0__n204), .C(
        n233), .Y(ALU_DW_rash_0__n743) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U312 ( .A(ALU_DW_rash_0__n77), .Y(ALU__N297) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U313 ( .A(ALU_DW_rash_0__n234), .Y(ALU_DW_rash_0__n233) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U314 ( .A(ALU_DW_rash_0__n625), .Y(ALU_DW_rash_0__n234) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U315 ( .A(ALU_DW_rash_0__n263), .Y(ALU_DW_rash_0__n235) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U316 ( .A(ALU_DW_rash_0__n237), .Y(ALU_DW_rash_0__n236) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U317 ( .A(ALU_DW_rash_0__n622), .Y(ALU_DW_rash_0__n237) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U318 ( .A(ALU_DW_rash_0__n239), .Y(ALU_DW_rash_0__n238) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U319 ( .A(ALU_DW_rash_0__n663), .Y(ALU_DW_rash_0__n239) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U320 ( .A(ALU_DW_rash_0__n655), .Y(ALU_DW_rash_0__n242) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U321 ( .A1(ALU_DW_rash_0__n310), .A2(ALU_DW_rash_0__n419), .B1(ALU_DW_rash_0__n255), .B2(ALU_DW_rash_0__n476), .Y(
        n651) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U322 ( .A(ALU_DW_rash_0__n123), .Y(ALU_DW_rash_0__n243) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U323 ( .A(ALU_DW_rash_0__n125), .Y(ALU_DW_rash_0__n244) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U324 ( .A1(ALU_DW_rash_0__n418), .A2(ALU_DW_rash_0__n433), .B1(ALU_DW_rash_0__n435), .B2(ALU_DW_rash_0__n204), .C(
        n246), .Y(ALU_DW_rash_0__n744) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U325 ( .A(ALU_DW_rash_0__n128), .Y(ALU__N296) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U326 ( .A(ALU_DW_rash_0__n247), .Y(ALU_DW_rash_0__n246) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U327 ( .A(ALU_DW_rash_0__n631), .Y(ALU_DW_rash_0__n247) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U328 ( .A(ALU_DW_rash_0__n720), .Y(ALU_DW_rash_0__n336) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U329 ( .A(ALU_DW_rash_0__n336), .Y(ALU__N322) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U330 ( .A(ALU_DW_rash_0__n250), .Y(ALU_DW_rash_0__n249) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U331 ( .A(ALU_DW_rash_0__n626), .Y(ALU_DW_rash_0__n250) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U332 ( .A(ALU_DW_rash_0__n252), .Y(ALU_DW_rash_0__n251) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U333 ( .A(ALU_DW_rash_0__n607), .Y(ALU_DW_rash_0__n252) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U334 ( .A(ALU_DW_rash_0__n251), .Y(ALU_DW_rash_0__n537) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U335 ( .A(ALU_DW_rash_0__n254), .Y(ALU_DW_rash_0__n253) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U336 ( .A(ALU_DW_rash_0__n68), .Y(ALU_DW_rash_0__n254) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U337 ( .A1(ALU_DW_rash_0__n424), .A2(ALU_DW_rash_0__n517), .B1(ALU_DW_rash_0__n462), .B2(ALU_DW_rash_0__n410), .C1(
        n376), .C2(ALU_DW_rash_0__n489), .Y(ALU_DW_rash_0__n653) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U338 ( .A(ALU_DW_rash_0__n61), .Y(ALU_DW_rash_0__n255) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U339 ( .A1(ALU_DW_rash_0__n390), .A2(ALU_DW_rash_0__n516), .B1(ALU_DW_rash_0__n326), .B2(ALU_DW_rash_0__n204), .C(
        n257), .Y(ALU_DW_rash_0__n745) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U340 ( .A(ALU_DW_rash_0__n135), .Y(ALU__N295) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U341 ( .A(ALU_DW_rash_0__n258), .Y(ALU_DW_rash_0__n257) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U342 ( .A(ALU_DW_rash_0__n634), .Y(ALU_DW_rash_0__n258) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U343 ( .A(ALU_DW_rash_0__n333), .Y(ALU_DW_rash_0__n259) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U344 ( .A(ALU_DW_rash_0__n333), .Y(ALU_DW_rash_0__n260) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U345 ( .A(ALU_DW_rash_0__n262), .Y(ALU_DW_rash_0__n261) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U346 ( .A(ALU_DW_rash_0__n600), .Y(ALU_DW_rash_0__n262) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U347 ( .A1(ALU_DW_rash_0__n553), .A2(ALU_DW_rash_0__n199), .B1(ALU_DW_rash_0__n565), .B2(ALU_DW_rash_0__n26), .C(
        n453), .Y(ALU_DW_rash_0__n600) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U348 ( .A(ALU_DW_rash_0__n266), .Y(ALU_DW_rash_0__n263) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U349 ( .A(ALU_DW_rash_0__n267), .Y(ALU_DW_rash_0__n264) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U350 ( .A(ALU_DW_rash_0__n268), .Y(ALU_DW_rash_0__n265) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U351 ( .A(ALU_DW_rash_0__n392), .Y(ALU_DW_rash_0__n266) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U352 ( .A(ALU_DW_rash_0__n392), .Y(ALU_DW_rash_0__n267) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U353 ( .A(ALU_DW_rash_0__n392), .Y(ALU_DW_rash_0__n268) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U354 ( .A(ALU__n969), .Y(ALU_DW_rash_0__n392) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U355 ( .A(ALU_DW_rash_0__n270), .Y(ALU_DW_rash_0__n269) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U356 ( .A(ALU_DW_rash_0__n121), .Y(ALU_DW_rash_0__n270) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U357 ( .A(ALU_DW_rash_0__n272), .Y(ALU_DW_rash_0__n271) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U358 ( .A(ALU_DW_rash_0__n657), .Y(ALU_DW_rash_0__n272) );
  AO22x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U359 ( .A1(ALU_DW_rash_0__n302), .A2(ALU_DW_rash_0__n580), .B1(ALU_DW_rash_0__n35), .B2(ALU_DW_rash_0__n589), .Y(ALU_DW_rash_0__n715) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U360 ( .A(ALU_DW_rash_0__n271), .Y(ALU_DW_rash_0__n509) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U361 ( .A1(ALU_DW_rash_0__n424), .A2(ALU_DW_rash_0__n461), .B1(ALU_DW_rash_0__n366), .B2(ALU_DW_rash_0__n203), .C(
        n274), .Y(ALU_DW_rash_0__n739) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U362 ( .A(ALU_DW_rash_0__n71), .Y(ALU__N301) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U363 ( .A(ALU_DW_rash_0__n275), .Y(ALU_DW_rash_0__n274) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U364 ( .A(ALU_DW_rash_0__n693), .Y(ALU_DW_rash_0__n275) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U365 ( .A(ALU_DW_rash_0__n729), .Y(ALU_DW_rash_0__n365) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U366 ( .A(ALU_DW_rash_0__n365), .Y(ALU__N311) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U367 ( .A(ALU_DW_rash_0__n726), .Y(ALU_DW_rash_0__n444) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U368 ( .A(ALU_DW_rash_0__n444), .Y(ALU__N314) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U369 ( .A(ALU__n731), .Y(ALU_DW_rash_0__n278) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U370 ( .A(ALU_DW_rash_0__n280), .Y(ALU_DW_rash_0__n279) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U371 ( .A(ALU_DW_rash_0__n611), .Y(ALU_DW_rash_0__n280) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U372 ( .A1(ALU_DW_rash_0__n298), .A2(ALU_DW_rash_0__n26), .B1(ALU_DW_rash_0__n569), .B2(n929), .C(
        n438), .Y(ALU_DW_rash_0__n611) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U373 ( .A(ALU_DW_rash_0__n282), .Y(ALU_DW_rash_0__n281) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U374 ( .A(ALU_DW_rash_0__n609), .Y(ALU_DW_rash_0__n282) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U375 ( .A(ALU_DW_rash_0__n284), .Y(ALU_DW_rash_0__n283) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U376 ( .A(ALU_DW_rash_0__n210), .Y(ALU_DW_rash_0__n284) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U377 ( .A(ALU_DW_rash_0__n286), .Y(ALU_DW_rash_0__n285) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U378 ( .A(ALU_DW_rash_0__n158), .Y(ALU_DW_rash_0__n286) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U379 ( .A1(ALU_DW_rash_0__n452), .A2(ALU_DW_rash_0__n517), .B1(ALU_DW_rash_0__n537), .B2(ALU_DW_rash_0__n410), .C1(
        n418), .C2(ALU_DW_rash_0__n163), .Y(ALU_DW_rash_0__n671) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U380 ( .A(ALU_DW_rash_0__n75), .Y(ALU_DW_rash_0__n287) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U381 ( .A1(ALU_DW_rash_0__n477), .A2(ALU_DW_rash_0__n307), .B1(ALU_DW_rash_0__n542), .B2(ALU_DW_rash_0__n147), .C(
        n289), .Y(ALU_DW_rash_0__n737) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U382 ( .A(ALU_DW_rash_0__n76), .Y(ALU__N303) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U383 ( .A(ALU_DW_rash_0__n290), .Y(ALU_DW_rash_0__n289) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U384 ( .A(ALU_DW_rash_0__n686), .Y(ALU_DW_rash_0__n290) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U385 ( .A(ALU_DW_rash_0__n534), .Y(ALU_DW_rash_0__n291) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U386 ( .A(ALU_DW_rash_0__n195), .Y(ALU_DW_rash_0__n292) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U387 ( .A(ALU_DW_rash_0__n194), .Y(ALU_DW_rash_0__n293) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U388 ( .A(ALU_DW_rash_0__n485), .Y(ALU_DW_rash_0__n294) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U389 ( .A(ALU_DW_rash_0__n296), .Y(ALU_DW_rash_0__n295) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U390 ( .A(ALU_DW_rash_0__n724), .Y(ALU_DW_rash_0__n296) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U391 ( .A(ALU_DW_rash_0__n298), .Y(ALU_DW_rash_0__n561) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U392 ( .A(ALU_DW_rash_0__n644), .Y(ALU_DW_rash_0__n298) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U393 ( .A(ALU_DW_rash_0__n337), .Y(ALU_DW_rash_0__n445) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U394 ( .A(ALU_DW_rash_0__n163), .Y(ALU_DW_rash_0__n488) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U395 ( .A(n1091), .Y(ALU_DW_rash_0__n299) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U396 ( .A(n1091), .Y(ALU_DW_rash_0__n300) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U397 ( .A(n1091), .Y(ALU_DW_rash_0__n301) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U398 ( .A(n1091), .Y(ALU_DW_rash_0__n302) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U399 ( .A(ALU_DW_rash_0__n179), .Y(ALU_DW_rash_0__n303) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U400 ( .A(ALU_DW_rash_0__n206), .Y(ALU_DW_rash_0__n306) );
  CKINVDCx14_ASAP7_75t_R ALU___ALU_DW_rash_0___U401 ( .A(ALU_DW_rash_0__n16), .Y(ALU_DW_rash_0__n549) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U402 ( .A(ALU_DW_rash_0__n49), .Y(ALU_DW_rash_0__n309) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U403 ( .A(ALU_DW_rash_0__n48), .Y(ALU_DW_rash_0__n311) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U404 ( .A(ALU_DW_rash_0__n727), .Y(ALU_DW_rash_0__n352) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U405 ( .A(ALU_DW_rash_0__n352), .Y(ALU__N313) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U406 ( .A(ALU__n794), .Y(ALU_DW_rash_0__n313) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U407 ( .A(ALU_DW_rash_0__n315), .Y(ALU_DW_rash_0__n314) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U408 ( .A(ALU_DW_rash_0__n261), .Y(ALU_DW_rash_0__n315) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U409 ( .A(ALU_DW_rash_0__n317), .Y(ALU_DW_rash_0__n316) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U410 ( .A(ALU_DW_rash_0__n616), .Y(ALU_DW_rash_0__n317) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U411 ( .A(ALU_DW_rash_0__n316), .Y(ALU_DW_rash_0__n493) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U412 ( .A(ALU_DW_rash_0__n319), .Y(ALU_DW_rash_0__n318) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U413 ( .A(ALU_DW_rash_0__n656), .Y(ALU_DW_rash_0__n319) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U414 ( .A1(ALU_DW_rash_0__n437), .A2(ALU_DW_rash_0__n517), .B1(ALU_DW_rash_0__n542), .B2(ALU_DW_rash_0__n410), .C1(
        n390), .C2(ALU_DW_rash_0__n489), .Y(ALU_DW_rash_0__n710) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U415 ( .A(ALU_DW_rash_0__n127), .Y(ALU_DW_rash_0__n320) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U416 ( .A1(ALU_DW_rash_0__n454), .A2(ALU_DW_rash_0__n549), .B1(ALU_DW_rash_0__n462), .B2(ALU_DW_rash_0__n147), .C(
        n322), .Y(ALU_DW_rash_0__n735) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U417 ( .A(ALU_DW_rash_0__n65), .Y(ALU__N305) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U418 ( .A(ALU_DW_rash_0__n323), .Y(ALU_DW_rash_0__n322) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U419 ( .A(ALU_DW_rash_0__n680), .Y(ALU_DW_rash_0__n323) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U420 ( .A(ALU_DW_rash_0__n730), .Y(ALU_DW_rash_0__n324) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U421 ( .A(ALU_DW_rash_0__n502), .Y(ALU__N310) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U422 ( .A(ALU_DW_rash_0__n329), .Y(ALU_DW_rash_0__n328) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U423 ( .A(ALU_DW_rash_0__n649), .Y(ALU_DW_rash_0__n329) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U424 ( .A(ALU_DW_rash_0__n328), .Y(ALU_DW_rash_0__n439) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U425 ( .A(ALU_DW_rash_0__n738), .Y(ALU_DW_rash_0__n330) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U426 ( .A(ALU_DW_rash_0__n347), .Y(ALU_DW_rash_0__n331) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U427 ( .A(ALU_DW_rash_0__n331), .Y(ALU_DW_rash_0__n594) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U428 ( .A(ALU_DW_rash_0__n425), .Y(ALU_DW_rash_0__n332) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U429 ( .A(ALU_DW_rash_0__n425), .Y(ALU_DW_rash_0__n333) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U430 ( .A(ALU_DW_rash_0__n425), .Y(ALU_DW_rash_0__n334) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U431 ( .A(ALU_DW_rash_0__n425), .Y(ALU_DW_rash_0__n335) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW_rash_0___U432 ( .A(ALU_DW_rash_0__n259), .B(ALU_DW_rash_0__n366), .Y(ALU__N317) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW_rash_0___U433 ( .A(ALU_DW_rash_0__n86), .B(ALU_DW_rash_0__n332), .Y(ALU__N316) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U434 ( .A(ALU_DW_rash_0__n148), .B(ALU_DW_rash_0__n492), .Y(ALU_DW_rash_0__n720) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U435 ( .A(ALU_DW_rash_0__n413), .Y(ALU_DW_rash_0__n337) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U436 ( .A(ALU_DW_rash_0__n339), .Y(ALU_DW_rash_0__n338) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U437 ( .A(ALU_DW_rash_0__n279), .Y(ALU_DW_rash_0__n339) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U438 ( .A(ALU_DW_rash_0__n160), .Y(ALU_DW_rash_0__n437) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U439 ( .A(n1010), .Y(ALU_DW_rash_0__n340) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U440 ( .A(n1010), .Y(ALU_DW_rash_0__n341) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U441 ( .A(ALU_DW_rash_0__n573), .Y(ALU_DW_rash_0__n567) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U442 ( .A(ALU_DW_rash_0__n200), .Y(ALU_DW_rash_0__n568) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U443 ( .A(ALU_DW_rash_0__n15), .Y(ALU_DW_rash_0__n569) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U444 ( .A(ALU_DW_rash_0__n575), .Y(ALU_DW_rash_0__n565) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U445 ( .A(ALU_DW_rash_0__n572), .Y(ALU_DW_rash_0__n566) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U446 ( .A(ALU_DW_rash_0__n303), .Y(ALU_DW_rash_0__n562) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U447 ( .A(n1174), .Y(ALU_DW_rash_0__n342) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW_rash_0___U448 ( .A(ALU_DW_rash_0__n344), .Y(ALU_DW_rash_0__n343) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U449 ( .A(ALU_DW_rash_0__n57), .Y(ALU_DW_rash_0__n344) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U450 ( .A1(ALU_DW_rash_0__n549), .A2(ALU_DW_rash_0__n440), .B1(ALU_DW_rash_0__n458), .B2(ALU_DW_rash_0__n393), .C(
        n346), .Y(ALU_DW_rash_0__n738) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U451 ( .A(ALU_DW_rash_0__n330), .Y(ALU__N302) );
  INVx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U452 ( .A(ALU_DW_rash_0__n594), .Y(ALU_DW_rash_0__n346) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U453 ( .A(ALU_DW_rash_0__n348), .Y(ALU_DW_rash_0__n347) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U454 ( .A(ALU_DW_rash_0__n1), .Y(ALU_DW_rash_0__n348) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U455 ( .A(ALU_DW_rash_0__n722), .Y(ALU_DW_rash_0__n501) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U456 ( .A(ALU_DW_rash_0__n501), .Y(ALU__N320) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U457 ( .A(ALU__n966), .Y(ALU_DW_rash_0__n389) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U458 ( .A(ALU_DW_rash_0__n728), .Y(ALU_DW_rash_0__n350) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U459 ( .A(ALU_DW_rash_0__n469), .Y(ALU__N312) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U460 ( .A(ALU_DW_rash_0__n240), .B(ALU_DW_rash_0__n334), .Y(ALU_DW_rash_0__n727) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U461 ( .A(ALU_DW_rash_0__n354), .Y(ALU_DW_rash_0__n353) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U462 ( .A(ALU_DW_rash_0__n660), .Y(ALU_DW_rash_0__n354) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U463 ( .A(ALU_DW_rash_0__n615), .Y(ALU_DW_rash_0__n355) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U464 ( .A1(ALU_DW_rash_0__n403), .A2(ALU_DW_rash_0__n549), .B1(ALU_DW_rash_0__n428), .B2(ALU_DW_rash_0__n458), .C(
        n504), .Y(ALU_DW_rash_0__n734) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U465 ( .A(ALU_DW_rash_0__n198), .Y(ALU_DW_rash_0__n356) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U466 ( .A(ALU_DW_rash_0__n358), .Y(ALU_DW_rash_0__n357) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U467 ( .A(ALU_DW_rash_0__n678), .Y(ALU_DW_rash_0__n358) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U468 ( .A(ALU_DW_rash_0__n357), .Y(ALU_DW_rash_0__n504) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U469 ( .A(ALU__n900), .Y(ALU_DW_rash_0__n359) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U470 ( .A(ALU__n900), .Y(ALU_DW_rash_0__n360) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U471 ( .A(ALU_DW_rash_0__n362), .Y(ALU_DW_rash_0__n361) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U472 ( .A(ALU_DW_rash_0__n645), .Y(ALU_DW_rash_0__n362) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U473 ( .A(ALU_DW_rash_0__n152), .Y(ALU_DW_rash_0__n363) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U474 ( .A(ALU_DW_rash_0__n725), .Y(ALU_DW_rash_0__n430) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U475 ( .A(ALU_DW_rash_0__n430), .Y(ALU__N315) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U476 ( .A(ALU_DW_rash_0__n326), .B(ALU_DW_rash_0__n260), .Y(ALU_DW_rash_0__n729) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U477 ( .A(ALU_DW_rash_0__n367), .Y(ALU_DW_rash_0__n366) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U478 ( .A(ALU_DW_rash_0__n353), .Y(ALU_DW_rash_0__n367) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U479 ( .A(ALU_DW_rash_0__n369), .Y(ALU_DW_rash_0__n368) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U480 ( .A(ALU_DW_rash_0__n605), .Y(ALU_DW_rash_0__n369) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U481 ( .A1(ALU_DW_rash_0__n363), .A2(ALU_DW_rash_0__n432), .B1(ALU_DW_rash_0__n269), .B2(ALU_DW_rash_0__n399), .C(
        n371), .Y(ALU_DW_rash_0__n742) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U482 ( .A(ALU_DW_rash_0__n107), .Y(ALU__N298) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U483 ( .A(ALU_DW_rash_0__n372), .Y(ALU_DW_rash_0__n371) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U484 ( .A(ALU_DW_rash_0__n619), .Y(ALU_DW_rash_0__n372) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U485 ( .A(ALU__n934), .Y(ALU_DW_rash_0__n373) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U486 ( .A(ALU_DW_rash_0__n375), .Y(ALU_DW_rash_0__n374) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U487 ( .A(ALU_DW_rash_0__n654), .Y(ALU_DW_rash_0__n375) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U488 ( .A(ALU_DW_rash_0__n311), .B(ALU_DW_rash_0__n58), .Y(ALU_DW_rash_0__n636) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U489 ( .A(ALU_DW_rash_0__n378), .Y(ALU_DW_rash_0__n377) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U490 ( .A(ALU_DW_rash_0__n395), .Y(ALU_DW_rash_0__n378) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U491 ( .A(ALU_DW_rash_0__n29), .Y(ALU_DW_rash_0__n381) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U492 ( .A(ALU_DW_rash_0__n30), .Y(ALU_DW_rash_0__n382) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U493 ( .A(ALU_DW_rash_0__n384), .Y(ALU_DW_rash_0__n383) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U494 ( .A(ALU_DW_rash_0__n83), .Y(ALU_DW_rash_0__n384) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U495 ( .A(n892), .B(ALU_DW_rash_0__n445), .Y(ALU_DW_rash_0__n547) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U496 ( .A(n1178), .Y(ALU_DW_rash_0__n385) );
  OR5x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U497 ( .A(ALU_DW_rash_0__n387), .B(n1162), .C(n1075), .D(n701), .E(
        n313), .Y(ALU_DW_rash_0__n703) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U498 ( .A(ALU_DW_rash_0__n81), .Y(ALU_DW_rash_0__n386) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U499 ( .A(ALU_DW_rash_0__n708), .Y(ALU_DW_rash_0__n387) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U500 ( .A(ALU__n966), .Y(ALU_DW_rash_0__n388) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U501 ( .A(ALU_DW_rash_0__n711), .Y(ALU_DW_rash_0__n391) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U502 ( .A(ALU_DW_rash_0__n691), .Y(ALU_DW_rash_0__n394) );
  CKINVDCx8_ASAP7_75t_R ALU___ALU_DW_rash_0___U503 ( .A(ALU_DW_rash_0__n526), .Y(ALU_DW_rash_0__n587) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U504 ( .A(ALU_DW_rash_0__n409), .Y(ALU_DW_rash_0__n395) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U505 ( .A(ALU_DW_rash_0__n377), .Y(ALU_DW_rash_0__n396) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U506 ( .A(ALU_DW_rash_0__n608), .Y(ALU_DW_rash_0__n397) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U507 ( .A(ALU_DW_rash_0__n399), .Y(ALU_DW_rash_0__n398) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U508 ( .A(ALU_DW_rash_0__n203), .Y(ALU_DW_rash_0__n399) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U509 ( .A1(ALU_DW_rash_0__n488), .A2(ALU_DW_rash_0__n464), .B1(ALU_DW_rash_0__n27), .B2(ALU_DW_rash_0__n493), .C(
        n401), .Y(ALU_DW_rash_0__n677) );
  INVx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U510 ( .A(ALU_DW_rash_0__n226), .Y(ALU_DW_rash_0__n400) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U511 ( .A(ALU_DW_rash_0__n402), .Y(ALU_DW_rash_0__n401) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U512 ( .A(ALU_DW_rash_0__n714), .Y(ALU_DW_rash_0__n402) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U513 ( .A(ALU_DW_rash_0__n690), .Y(ALU_DW_rash_0__n404) );
  CKINVDCx8_ASAP7_75t_R ALU___ALU_DW_rash_0___U514 ( .A(ALU_DW_rash_0__n585), .Y(ALU_DW_rash_0__n536) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U515 ( .A(ALU_DW_rash_0__n482), .Y(ALU_DW_rash_0__n521) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U516 ( .A(ALU_DW_rash_0__n548), .B(ALU_DW_rash_0__n379), .Y(ALU_DW_rash_0__n694) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U517 ( .A(ALU__n1032), .Y(ALU_DW_rash_0__n405) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U518 ( .A(ALU__n1032), .Y(ALU_DW_rash_0__n406) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U519 ( .A(ALU__n1035), .Y(ALU_DW_rash_0__n407) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U520 ( .A(ALU_DW_rash_0__n396), .Y(ALU_DW_rash_0__n408) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U521 ( .A(ALU_DW_rash_0__n397), .Y(ALU_DW_rash_0__n409) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U522 ( .A(ALU_DW_rash_0__n359), .B(ALU_DW_rash_0__n264), .Y(ALU_DW_rash_0__n642) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U523 ( .A(ALU_DW_rash_0__n723), .Y(ALU_DW_rash_0__n411) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U524 ( .A(ALU_DW_rash_0__n540), .Y(ALU__N319) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U525 ( .A(ALU_DW_rash_0__n596), .Y(ALU_DW_rash_0__n413) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U526 ( .A(ALU_DW_rash_0__n415), .Y(ALU_DW_rash_0__n414) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U527 ( .A(ALU_DW_rash_0__n661), .Y(ALU_DW_rash_0__n415) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U528 ( .A(ALU_DW_rash_0__n417), .Y(ALU_DW_rash_0__n416) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U529 ( .A(ALU_DW_rash_0__n672), .Y(ALU_DW_rash_0__n417) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U530 ( .A1(ALU_DW_rash_0__n410), .A2(ALU_DW_rash_0__n439), .B1(ALU_DW_rash_0__n517), .B2(ALU_DW_rash_0__n454), .C(
        n420), .Y(ALU_DW_rash_0__n652) );
  INVx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U531 ( .A(ALU_DW_rash_0__n138), .Y(ALU_DW_rash_0__n419) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U532 ( .A(ALU_DW_rash_0__n421), .Y(ALU_DW_rash_0__n420) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U533 ( .A(ALU_DW_rash_0__n675), .Y(ALU_DW_rash_0__n421) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U534 ( .A(ALU_DW_rash_0__n423), .Y(ALU_DW_rash_0__n422) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U535 ( .A(ALU_DW_rash_0__n699), .Y(ALU_DW_rash_0__n423) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U536 ( .A(ALU_DW_rash_0__n379), .Y(ALU_DW_rash_0__n425) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U537 ( .A(ALU_DW_rash_0__n427), .Y(ALU_DW_rash_0__n426) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U538 ( .A(ALU_DW_rash_0__n658), .Y(ALU_DW_rash_0__n427) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U539 ( .A1(n1182), .A2(ALU_DW_rash_0__n577), .B1(ALU_DW_rash_0__n388), .B2(ALU_DW_rash_0__n585), .C(
        n429), .Y(ALU_DW_rash_0__n622) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U540 ( .A(ALU_DW_rash_0__n689), .Y(ALU_DW_rash_0__n429) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U541 ( .A(ALU_DW_rash_0__n154), .B(ALU_DW_rash_0__n381), .Y(ALU_DW_rash_0__n725) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U542 ( .A(ALU_DW_rash_0__n647), .Y(ALU_DW_rash_0__n431) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U543 ( .A(ALU_DW_rash_0__n460), .Y(ALU_DW_rash_0__n432) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U544 ( .A(ALU_DW_rash_0__n460), .Y(ALU_DW_rash_0__n433) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW_rash_0___U545 ( .A(n1114), .Y(ALU_DW_rash_0__n434) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U546 ( .A(ALU_DW_rash_0__n713), .Y(ALU_DW_rash_0__n438) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U547 ( .A1(ALU_DW_rash_0__n472), .A2(ALU_DW_rash_0__n577), .B1(ALU_DW_rash_0__n199), .B2(ALU_DW_rash_0__n586), .Y(
        n713) );
  AO22x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U548 ( .A1(ALU_DW_rash_0__n562), .A2(ALU_DW_rash_0__n340), .B1(ALU_DW_rash_0__n550), .B2(ALU_DW_rash_0__n300), .Y(
        n649) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U549 ( .A1(ALU_DW_rash_0__n551), .A2(n1064), .B1(ALU_DW_rash_0__n564), .B2(ALU_DW_rash_0__n385), .C(
        n441), .Y(ALU_DW_rash_0__n665) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U550 ( .A(ALU_DW_rash_0__n692), .Y(ALU_DW_rash_0__n441) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U551 ( .A(ALU_DW_rash_0__n443), .Y(ALU_DW_rash_0__n442) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U552 ( .A(ALU_DW_rash_0__n721), .Y(ALU_DW_rash_0__n443) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U553 ( .A(ALU_DW_rash_0__n269), .B(ALU_DW_rash_0__n382), .Y(ALU_DW_rash_0__n726) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U554 ( .A(n749), .Y(ALU_DW_rash_0__n596) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U555 ( .A1(ALU_DW_rash_0__n437), .A2(ALU_DW_rash_0__n459), .B1(ALU_DW_rash_0__n154), .B2(ALU_DW_rash_0__n167), .C(
        n447), .Y(ALU_DW_rash_0__n741) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U556 ( .A(ALU_DW_rash_0__n89), .Y(ALU__N299) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U557 ( .A(ALU_DW_rash_0__n448), .Y(ALU_DW_rash_0__n447) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U558 ( .A(ALU_DW_rash_0__n613), .Y(ALU_DW_rash_0__n448) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U559 ( .A1(ALU_DW_rash_0__n410), .A2(ALU_DW_rash_0__n544), .B1(ALU_DW_rash_0__n517), .B2(ALU_DW_rash_0__n466), .C(
        n450), .Y(ALU_DW_rash_0__n670) );
  INVx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U560 ( .A(ALU_DW_rash_0__n208), .Y(ALU_DW_rash_0__n449) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U561 ( .A(ALU_DW_rash_0__n451), .Y(ALU_DW_rash_0__n450) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U562 ( .A(ALU_DW_rash_0__n676), .Y(ALU_DW_rash_0__n451) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U563 ( .A(ALU_DW_rash_0__n673), .Y(ALU_DW_rash_0__n453) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U564 ( .A1(ALU_DW_rash_0__n553), .A2(n1160), .B1(ALU_DW_rash_0__n567), .B2(n1100), .C(
        n455), .Y(ALU_DW_rash_0__n666) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U565 ( .A(ALU_DW_rash_0__n698), .Y(ALU_DW_rash_0__n455) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U566 ( .A1(ALU_DW_rash_0__n550), .A2(n1068), .B1(ALU_DW_rash_0__n570), .B2(ALU_DW_rash_0__n407), .C(
        n457), .Y(ALU_DW_rash_0__n620) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U567 ( .A(ALU_DW_rash_0__n688), .Y(ALU_DW_rash_0__n457) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U568 ( .A(ALU_DW_rash_0__n433), .Y(ALU_DW_rash_0__n458) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U569 ( .A(ALU_DW_rash_0__n432), .Y(ALU_DW_rash_0__n459) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U570 ( .A(ALU_DW_rash_0__n516), .Y(ALU_DW_rash_0__n460) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U571 ( .A(ALU_DW_rash_0__n601), .Y(ALU_DW_rash_0__n461) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U572 ( .A1(ALU_DW_rash_0__n389), .A2(ALU_DW_rash_0__n577), .B1(ALU_DW_rash_0__n585), .B2(ALU_DW_rash_0__n150), .C(
        n463), .Y(ALU_DW_rash_0__n628) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U573 ( .A(ALU_DW_rash_0__n696), .Y(ALU_DW_rash_0__n463) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U574 ( .A1(ALU_DW_rash_0__n555), .A2(n1225), .B1(ALU_DW_rash_0__n569), .B2(n1068), .C(
        n465), .Y(ALU_DW_rash_0__n614) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U575 ( .A(ALU_DW_rash_0__n718), .Y(ALU_DW_rash_0__n465) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U576 ( .A1(ALU_DW_rash_0__n552), .A2(n1100), .B1(ALU_DW_rash_0__n566), .B2(ALU_DW_rash_0__n373), .C(
        n467), .Y(ALU_DW_rash_0__n661) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U577 ( .A(ALU_DW_rash_0__n685), .Y(ALU_DW_rash_0__n467) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U578 ( .A(ALU_DW_rash_0__n732), .Y(ALU__N308) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U579 ( .A(ALU_DW_rash_0__n435), .B(ALU_DW_rash_0__n380), .Y(ALU_DW_rash_0__n728) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U580 ( .A(ALU_DW_rash_0__n350), .Y(ALU_DW_rash_0__n469) );
  O2A1O1Ixp33_ASAP7_75t_R ALU___ALU_DW_rash_0___U581 ( .A1(ALU_DW_rash_0__n212), .A2(ALU_DW_rash_0__n172), .B(ALU_DW_rash_0__n213), .C(ALU_DW_rash_0__n497), .Y(
        N291) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U582 ( .A(n1152), .Y(ALU_DW_rash_0__n470) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U583 ( .A(n1152), .Y(ALU_DW_rash_0__n471) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U584 ( .A(n1152), .Y(ALU_DW_rash_0__n472) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U585 ( .A1(ALU_DW_rash_0__n466), .A2(ALU_DW_rash_0__n549), .B1(ALU_DW_rash_0__n537), .B2(ALU_DW_rash_0__n148), .C(
        n474), .Y(ALU_DW_rash_0__n736) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U586 ( .A(ALU_DW_rash_0__n120), .Y(ALU__N304) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U587 ( .A(ALU_DW_rash_0__n475), .Y(ALU_DW_rash_0__n474) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U588 ( .A(ALU_DW_rash_0__n681), .Y(ALU_DW_rash_0__n475) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U589 ( .A(ALU_DW_rash_0__n359), .Y(ALU_DW_rash_0__n598) );
  CKINVDCx5p33_ASAP7_75t_R ALU___ALU_DW_rash_0___U590 ( .A(ALU_DW_rash_0__n599), .Y(ALU_DW_rash_0__n476) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U591 ( .A1(ALU_DW_rash_0__n553), .A2(ALU_DW_rash_0__n373), .B1(ALU_DW_rash_0__n569), .B2(n1064), .C(
        n478), .Y(ALU_DW_rash_0__n663) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U592 ( .A(ALU_DW_rash_0__n716), .Y(ALU_DW_rash_0__n478) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U593 ( .A1(ALU_DW_rash_0__n552), .A2(ALU_DW_rash_0__n407), .B1(ALU_DW_rash_0__n563), .B2(n1182), .C(
        n480), .Y(ALU_DW_rash_0__n626) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U594 ( .A(ALU_DW_rash_0__n249), .Y(ALU_DW_rash_0__n479) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U595 ( .A(ALU_DW_rash_0__n695), .Y(ALU_DW_rash_0__n480) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U596 ( .A(ALU_DW_rash_0__n482), .Y(ALU_DW_rash_0__n481) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U597 ( .A(ALU_DW_rash_0__n483), .Y(ALU_DW_rash_0__n482) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U598 ( .A(ALU_DW_rash_0__n524), .Y(ALU_DW_rash_0__n483) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U599 ( .A(ALU_DW_rash_0__n556), .Y(ALU_DW_rash_0__n524) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U600 ( .A(ALU_DW_rash_0__n51), .Y(ALU_DW_rash_0__n484) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U601 ( .A(ALU_DW_rash_0__n545), .Y(ALU_DW_rash_0__n485) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U602 ( .A(ALU_DW_rash_0__n584), .Y(ALU_DW_rash_0__n583) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U603 ( .A(ALU_DW_rash_0__n484), .Y(ALU_DW_rash_0__n545) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U604 ( .A(ALU_DW_rash_0__n694), .Y(ALU_DW_rash_0__n486) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U605 ( .A(ALU_DW_rash_0__n679), .Y(ALU_DW_rash_0__n487) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U606 ( .A(n892), .B(n749), .Y(ALU_DW_rash_0__n646) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U607 ( .A(ALU_DW_rash_0__n445), .B(n892), .Y(ALU_DW_rash_0__n644) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U608 ( .A(ALU_DW_rash_0__n164), .Y(ALU_DW_rash_0__n489) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U609 ( .A(ALU_DW_rash_0__n731), .Y(ALU__N309) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U610 ( .A(ALU_DW_rash_0__n299), .B(ALU_DW_rash_0__n562), .Y(ALU_DW_rash_0__n648) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U611 ( .A1(ALU_DW_rash_0__n555), .A2(ALU_DW_rash_0__n389), .B1(ALU_DW_rash_0__n150), .B2(ALU_DW_rash_0__n570), .C(
        n494), .Y(ALU_DW_rash_0__n616) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U612 ( .A(ALU_DW_rash_0__n717), .Y(ALU_DW_rash_0__n494) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U613 ( .A1(ALU_DW_rash_0__n550), .A2(n1024), .B1(ALU_DW_rash_0__n565), .B2(n1225), .C(
        n496), .Y(ALU_DW_rash_0__n605) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U614 ( .A(ALU_DW_rash_0__n683), .Y(ALU_DW_rash_0__n496) );
  AND4x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U615 ( .A(ALU_DW_rash_0__n188), .B(ALU_DW_rash_0__n386), .C(ALU_DW_rash_0__n499), .D(ALU_DW_rash_0__n500), .Y(ALU_DW_rash_0__n638)
         );
  OR4x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U616 ( .A(ALU_DW_rash_0__n12), .B(n1164), .C(n352), .D(ALU_DW_rash_0__n20), .Y(ALU_DW_rash_0__n702)
         );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U617 ( .A(ALU_DW_rash_0__n186), .Y(ALU_DW_rash_0__n498) );
  OR5x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U618 ( .A(ALU_DW_rash_0__n10), .B(n1123), .C(n1033), .D(ALU_DW_rash_0__n93), .E(n978), .Y(ALU_DW_rash_0__n704) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U619 ( .A(ALU_DW_rash_0__n189), .Y(ALU_DW_rash_0__n499) );
  OR5x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U620 ( .A(ALU_DW_rash_0__n11), .B(n1208), .C(n619), .D(ALU_DW_rash_0__n67), .E(ALU_DW_rash_0__n13), 
        .Y(ALU_DW_rash_0__n705) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U621 ( .A(ALU_DW_rash_0__n191), .Y(ALU_DW_rash_0__n500) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U622 ( .A(ALU_DW_rash_0__n544), .B(ALU_DW_rash_0__n149), .Y(ALU_DW_rash_0__n722) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U623 ( .A(ALU_DW_rash_0__n253), .B(ALU_DW_rash_0__n381), .Y(ALU_DW_rash_0__n730) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U624 ( .A(ALU_DW_rash_0__n324), .Y(ALU_DW_rash_0__n502) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U625 ( .A(ALU_DW_rash_0__n356), .Y(ALU__N306) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U626 ( .A1(ALU_DW_rash_0__n552), .A2(n1182), .B1(ALU_DW_rash_0__n563), .B2(ALU_DW_rash_0__n388), .C(
        n506), .Y(ALU_DW_rash_0__n609) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U627 ( .A(ALU_DW_rash_0__n682), .Y(ALU_DW_rash_0__n506) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U628 ( .A1(ALU_DW_rash_0__n553), .A2(ALU_DW_rash_0__n385), .B1(ALU_DW_rash_0__n562), .B2(n1024), .C(
        n508), .Y(ALU_DW_rash_0__n667) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U629 ( .A(ALU_DW_rash_0__n697), .Y(ALU_DW_rash_0__n508) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U630 ( .A1(ALU_DW_rash_0__n551), .A2(n1215), .B1(ALU_DW_rash_0__n566), .B2(n920), .C(
        n510), .Y(ALU_DW_rash_0__n657) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U631 ( .A(ALU_DW_rash_0__n715), .Y(ALU_DW_rash_0__n510) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW_rash_0___U632 ( .A(ALU_DW_rash_0__n527), .Y(ALU_DW_rash_0__n511) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U633 ( .A(ALU_DW_rash_0__n530), .Y(ALU_DW_rash_0__n527) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U634 ( .A(ALU_DW_rash_0__n581), .Y(ALU_DW_rash_0__n512) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U635 ( .A(ALU_DW_rash_0__n582), .Y(ALU_DW_rash_0__n513) );
  CKINVDCx5p33_ASAP7_75t_R ALU___ALU_DW_rash_0___U636 ( .A(ALU_DW_rash_0__n513), .Y(ALU_DW_rash_0__n577) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U637 ( .A(ALU_DW_rash_0__n292), .Y(ALU_DW_rash_0__n581) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U638 ( .A(ALU_DW_rash_0__n560), .Y(ALU_DW_rash_0__n558) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U639 ( .A(n749), .B(n892), .Y(ALU_DW_rash_0__n514) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U640 ( .A(ALU_DW_rash_0__n459), .Y(ALU_DW_rash_0__n515) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U641 ( .A(ALU_DW_rash_0__n461), .Y(ALU_DW_rash_0__n516) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U642 ( .A(ALU_DW_rash_0__n360), .B(ALU_DW_rash_0__n597), .Y(ALU_DW_rash_0__n641) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U643 ( .A(ALU_DW_rash_0__n733), .Y(ALU__N307) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U644 ( .A(ALU_DW_rash_0__n439), .B(ALU_DW_rash_0__n148), .Y(ALU_DW_rash_0__n721) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U645 ( .A(ALU_DW_rash_0__n442), .Y(ALU__N321) );
  OR3x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U646 ( .A(ALU_DW_rash_0__n381), .B(ALU_DW_rash_0__n360), .C(ALU_DW_rash_0__n285), .Y(ALU_DW_rash_0__n724) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U647 ( .A(ALU_DW_rash_0__n295), .Y(ALU__N318) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U648 ( .A(ALU_DW_rash_0__n581), .Y(ALU_DW_rash_0__n579) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U649 ( .A(ALU_DW_rash_0__n293), .Y(ALU_DW_rash_0__n582) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U650 ( .A(ALU_DW_rash_0__n512), .Y(ALU_DW_rash_0__n578) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U651 ( .A(ALU_DW_rash_0__n175), .Y(ALU_DW_rash_0__n522) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U652 ( .A(ALU_DW_rash_0__n175), .Y(ALU_DW_rash_0__n523) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U653 ( .A(ALU_DW_rash_0__n197), .Y(ALU_DW_rash_0__n525) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U654 ( .A(ALU_DW_rash_0__n99), .Y(ALU_DW_rash_0__n556) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U655 ( .A(ALU_DW_rash_0__n536), .Y(ALU_DW_rash_0__n528) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U656 ( .A(ALU_DW_rash_0__n174), .Y(ALU_DW_rash_0__n529) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U657 ( .A(ALU_DW_rash_0__n173), .Y(ALU_DW_rash_0__n530) );
  INVx5_ASAP7_75t_R ALU___ALU_DW_rash_0___U658 ( .A(ALU_DW_rash_0__n528), .Y(ALU_DW_rash_0__n586) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U659 ( .A(ALU_DW_rash_0__n593), .Y(ALU_DW_rash_0__n592) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U660 ( .A(ALU_DW_rash_0__n486), .B(ALU_DW_rash_0__n597), .Y(ALU_DW_rash_0__n610) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW_rash_0___U661 ( .A(ALU_DW_rash_0__n533), .Y(ALU_DW_rash_0__n532) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW_rash_0___U662 ( .A(ALU_DW_rash_0__n595), .Y(ALU_DW_rash_0__n533) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U663 ( .A(ALU_DW_rash_0__n536), .Y(ALU_DW_rash_0__n534) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U664 ( .A(ALU_DW_rash_0__n591), .Y(ALU_DW_rash_0__n535) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U665 ( .A(ALU_DW_rash_0__n291), .Y(ALU_DW_rash_0__n588) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U666 ( .A(ALU_DW_rash_0__n546), .Y(ALU_DW_rash_0__n591) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U667 ( .A(ALU_DW_rash_0__n557), .Y(ALU_DW_rash_0__n551) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U668 ( .A(ALU_DW_rash_0__n100), .Y(ALU_DW_rash_0__n557) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U669 ( .A1(ALU_DW_rash_0__n555), .A2(n969), .B1(ALU_DW_rash_0__n564), .B2(ALU_DW_rash_0__n38), .C(
        n538), .Y(ALU_DW_rash_0__n607) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U670 ( .A(ALU_DW_rash_0__n684), .Y(ALU_DW_rash_0__n538) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U671 ( .A(ALU_DW_rash_0__n548), .B(ALU_DW_rash_0__n597), .Y(ALU_DW_rash_0__n662) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U672 ( .A(ALU_DW_rash_0__n509), .B(ALU_DW_rash_0__n149), .Y(ALU_DW_rash_0__n723) );
  INVx1_ASAP7_75t_R ALU___ALU_DW_rash_0___U673 ( .A(ALU_DW_rash_0__n411), .Y(ALU_DW_rash_0__n540) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U674 ( .A(ALU_DW_rash_0__n382), .Y(ALU_DW_rash_0__n595) );
  INVx3_ASAP7_75t_R ALU___ALU_DW_rash_0___U675 ( .A(ALU_DW_rash_0__n532), .Y(ALU_DW_rash_0__n541) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U676 ( .A1(ALU_DW_rash_0__n552), .A2(ALU_DW_rash_0__n38), .B1(ALU_DW_rash_0__n568), .B2(n1109), .C(
        n543), .Y(ALU_DW_rash_0__n615) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW_rash_0___U677 ( .A(ALU_DW_rash_0__n712), .Y(ALU_DW_rash_0__n543) );
  AO222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U678 ( .A1(ALU_DW_rash_0__n550), .A2(ALU_DW_rash_0__n340), .B1(ALU_DW_rash_0__n586), .B2(ALU_DW_rash_0__n301), .C1(
        n562), .C2(n1215), .Y(ALU_DW_rash_0__n656) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U679 ( .A(ALU_DW_rash_0__n318), .Y(ALU_DW_rash_0__n544) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U680 ( .A(ALU_DW_rash_0__n559), .Y(ALU_DW_rash_0__n555) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U681 ( .A(ALU_DW_rash_0__n560), .Y(ALU_DW_rash_0__n559) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U682 ( .A(ALU_DW_rash_0__n297), .Y(ALU_DW_rash_0__n560) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U683 ( .A(ALU_DW_rash_0__n523), .Y(ALU_DW_rash_0__n553) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U684 ( .A(ALU_DW_rash_0__n14), .Y(ALU_DW_rash_0__n570) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U685 ( .A(ALU_DW_rash_0__n22), .Y(ALU_DW_rash_0__n571) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U686 ( .A(ALU_DW_rash_0__n104), .Y(ALU_DW_rash_0__n576) );
  INVx4_ASAP7_75t_R ALU___ALU_DW_rash_0___U687 ( .A(ALU_DW_rash_0__n587), .Y(ALU_DW_rash_0__n546) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW_rash_0___U688 ( .A(ALU_DW_rash_0__n547), .Y(ALU_DW_rash_0__n593) );
  INVx6_ASAP7_75t_R ALU___ALU_DW_rash_0___U689 ( .A(ALU_DW_rash_0__n598), .Y(ALU_DW_rash_0__n548) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U690 ( .A(ALU_DW_rash_0__n486), .B(ALU_DW_rash_0__n265), .Y(ALU_DW_rash_0__n606) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW_rash_0___U691 ( .A(ALU_DW_rash_0__n335), .B(ALU_DW_rash_0__n488), .Y(ALU_DW_rash_0__n608) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U692 ( .A1(ALU_DW_rash_0__n495), .A2(ALU_DW_rash_0__n549), .B1(ALU_DW_rash_0__n537), .B2(ALU_DW_rash_0__n409), .C1(
        n505), .C2(ALU_DW_rash_0__n182), .Y(ALU_DW_rash_0__n604) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U693 ( .A1(ALU_DW_rash_0__n464), .A2(ALU_DW_rash_0__n549), .B1(ALU_DW_rash_0__n542), .B2(ALU_DW_rash_0__n378), .C1(
        n493), .C2(ALU_DW_rash_0__n183), .Y(ALU_DW_rash_0__n613) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U694 ( .A1(ALU_DW_rash_0__n456), .A2(ALU_DW_rash_0__n549), .B1(ALU_DW_rash_0__n393), .B2(ALU_DW_rash_0__n396), .C1(
        n428), .C2(ALU_DW_rash_0__n182), .Y(ALU_DW_rash_0__n619) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U695 ( .A1(ALU_DW_rash_0__n479), .A2(ALU_DW_rash_0__n549), .B1(ALU_DW_rash_0__n424), .B2(ALU_DW_rash_0__n397), .C1(
        n462), .C2(ALU_DW_rash_0__n183), .Y(ALU_DW_rash_0__n625) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U696 ( .A1(ALU_DW_rash_0__n505), .A2(ALU_DW_rash_0__n549), .B1(ALU_DW_rash_0__n452), .B2(ALU_DW_rash_0__n377), .C1(
        n537), .C2(ALU_DW_rash_0__n183), .Y(ALU_DW_rash_0__n631) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U697 ( .A1(ALU_DW_rash_0__n493), .A2(ALU_DW_rash_0__n307), .B1(ALU_DW_rash_0__n437), .B2(ALU_DW_rash_0__n408), .C1(
        n542), .C2(ALU_DW_rash_0__n183), .Y(ALU_DW_rash_0__n634) );
  O2A1O1Ixp33_ASAP7_75t_R ALU___ALU_DW_rash_0___U698 ( .A1(ALU_DW_rash_0__n221), .A2(ALU_DW_rash_0__n172), .B(ALU_DW_rash_0__n219), .C(ALU_DW_rash_0__n497), .Y(
        N294) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U699 ( .A1(ALU_DW_rash_0__n476), .A2(ALU_DW_rash_0__n253), .B1(ALU_DW_rash_0__n220), .B2(ALU_DW_rash_0__n309), .Y(
        n637) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U700 ( .A1(ALU_DW_rash_0__n393), .A2(ALU_DW_rash_0__n517), .B1(ALU_DW_rash_0__n428), .B2(ALU_DW_rash_0__n410), .C1(
        n363), .C2(ALU_DW_rash_0__n106), .Y(ALU_DW_rash_0__n640) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U701 ( .A1(ALU_DW_rash_0__n199), .A2(ALU_DW_rash_0__n177), .B1(ALU_DW_rash_0__n26), .B2(ALU_DW_rash_0__n590), .Y(ALU_DW_rash_0__n645) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U702 ( .A1(ALU_DW_rash_0__n590), .A2(n1233), .B1(ALU_DW_rash_0__n578), .B2(n973), .Y(
        n647) );
  O2A1O1Ixp33_ASAP7_75t_R ALU___ALU_DW_rash_0___U703 ( .A1(ALU_DW_rash_0__n244), .A2(ALU_DW_rash_0__n172), .B(ALU_DW_rash_0__n243), .C(ALU_DW_rash_0__n497), .Y(
        N293) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U704 ( .A1(ALU_DW_rash_0__n26), .A2(ALU_DW_rash_0__n579), .B1(n929), .B2(ALU_DW_rash_0__n586), .Y(ALU_DW_rash_0__n654) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U705 ( .A1(ALU_DW_rash_0__n590), .A2(ALU_DW_rash_0__n342), .B1(ALU_DW_rash_0__n578), .B2(n1233), .Y(
        n655) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U706 ( .A1(ALU_DW_rash_0__n466), .A2(ALU_DW_rash_0__n59), .B1(ALU_DW_rash_0__n544), .B2(ALU_DW_rash_0__n489), .Y(ALU_DW_rash_0__n602) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U707 ( .A1(ALU_DW_rash_0__n477), .A2(ALU_DW_rash_0__n60), .B1(ALU_DW_rash_0__n509), .B2(ALU_DW_rash_0__n105), .Y(ALU_DW_rash_0__n612) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U708 ( .A1(ALU_DW_rash_0__n403), .A2(ALU_DW_rash_0__n162), .B1(ALU_DW_rash_0__n492), .B2(ALU_DW_rash_0__n517), .C1(
        n440), .C2(ALU_DW_rash_0__n60), .Y(ALU_DW_rash_0__n618) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U709 ( .A1(ALU_DW_rash_0__n454), .A2(ALU_DW_rash_0__n489), .B1(ALU_DW_rash_0__n439), .B2(ALU_DW_rash_0__n517), .C1(
        n507), .C2(ALU_DW_rash_0__n60), .Y(ALU_DW_rash_0__n624) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U710 ( .A1(ALU_DW_rash_0__n466), .A2(ALU_DW_rash_0__n488), .B1(ALU_DW_rash_0__n544), .B2(ALU_DW_rash_0__n517), .C1(
        n495), .C2(ALU_DW_rash_0__n59), .Y(ALU_DW_rash_0__n630) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U711 ( .A1(ALU_DW_rash_0__n477), .A2(ALU_DW_rash_0__n488), .B1(ALU_DW_rash_0__n509), .B2(ALU_DW_rash_0__n517), .C1(
        n464), .C2(ALU_DW_rash_0__n59), .Y(ALU_DW_rash_0__n633) );
  O2A1O1Ixp33_ASAP7_75t_R ALU___ALU_DW_rash_0___U712 ( .A1(ALU_DW_rash_0__n231), .A2(ALU_DW_rash_0__n172), .B(ALU_DW_rash_0__n230), .C(ALU_DW_rash_0__n497), .Y(
        N292) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U713 ( .A1(n929), .A2(ALU_DW_rash_0__n579), .B1(ALU_DW_rash_0__n434), .B2(ALU_DW_rash_0__n586), .Y(
        n672) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U714 ( .A1(n1109), .A2(ALU_DW_rash_0__n579), .B1(ALU_DW_rash_0__n471), .B2(ALU_DW_rash_0__n586), .Y(
        n673) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U715 ( .A1(ALU_DW_rash_0__n590), .A2(n1060), .B1(ALU_DW_rash_0__n578), .B2(ALU_DW_rash_0__n342), .Y(
        n674) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U716 ( .A1(ALU_DW_rash_0__n60), .A2(ALU_DW_rash_0__n456), .B1(ALU_DW_rash_0__n164), .B2(ALU_DW_rash_0__n440), .C1(
        n548), .C2(ALU_DW_rash_0__n285), .Y(ALU_DW_rash_0__n639) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U717 ( .A(ALU_DW_rash_0__n419), .B(ALU_DW_rash_0__n541), .Y(ALU_DW_rash_0__n731) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U718 ( .A1(ALU_DW_rash_0__n479), .A2(ALU_DW_rash_0__n60), .B1(ALU_DW_rash_0__n507), .B2(ALU_DW_rash_0__n166), .Y(ALU_DW_rash_0__n675) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U719 ( .A(ALU_DW_rash_0__n449), .B(ALU_DW_rash_0__n541), .Y(ALU_DW_rash_0__n732) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U720 ( .A1(ALU_DW_rash_0__n505), .A2(ALU_DW_rash_0__n59), .B1(ALU_DW_rash_0__n495), .B2(ALU_DW_rash_0__n489), .Y(ALU_DW_rash_0__n676) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U721 ( .A(ALU_DW_rash_0__n400), .B(ALU_DW_rash_0__n541), .Y(ALU_DW_rash_0__n733) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U722 ( .A1(ALU_DW_rash_0__n182), .A2(ALU_DW_rash_0__n440), .B1(ALU_DW_rash_0__n487), .B2(ALU_DW_rash_0__n492), .C1(
        n408), .C2(ALU_DW_rash_0__n456), .Y(ALU_DW_rash_0__n678) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U723 ( .A1(ALU_DW_rash_0__n182), .A2(ALU_DW_rash_0__n507), .B1(ALU_DW_rash_0__n487), .B2(ALU_DW_rash_0__n439), .C1(
        n408), .C2(ALU_DW_rash_0__n479), .Y(ALU_DW_rash_0__n680) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U724 ( .A1(ALU_DW_rash_0__n182), .A2(ALU_DW_rash_0__n495), .B1(ALU_DW_rash_0__n487), .B2(ALU_DW_rash_0__n544), .C1(
        n408), .C2(ALU_DW_rash_0__n505), .Y(ALU_DW_rash_0__n681) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U725 ( .A1(n1068), .A2(ALU_DW_rash_0__n578), .B1(ALU_DW_rash_0__n407), .B2(ALU_DW_rash_0__n586), .Y(
        n682) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U726 ( .A1(n1064), .A2(ALU_DW_rash_0__n580), .B1(ALU_DW_rash_0__n385), .B2(ALU_DW_rash_0__n588), .Y(
        n683) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U727 ( .A1(ALU_DW_rash_0__n150), .A2(ALU_DW_rash_0__n580), .B1(n925), .B2(ALU_DW_rash_0__n589), .Y(
        n684) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U728 ( .A1(n920), .A2(ALU_DW_rash_0__n177), .B1(n1160), .B2(ALU_DW_rash_0__n590), .Y(
        n685) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U729 ( .A1(ALU_DW_rash_0__n182), .A2(ALU_DW_rash_0__n464), .B1(ALU_DW_rash_0__n487), .B2(ALU_DW_rash_0__n509), .C1(
        n408), .C2(ALU_DW_rash_0__n493), .Y(ALU_DW_rash_0__n686) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U730 ( .A1(n1024), .A2(ALU_DW_rash_0__n72), .B1(n1225), .B2(ALU_DW_rash_0__n587), .Y(
        n688) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U731 ( .A1(n925), .A2(ALU_DW_rash_0__n563), .B1(ALU_DW_rash_0__n150), .B2(ALU_DW_rash_0__n554), .Y(
        n689) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U732 ( .A1(ALU_DW_rash_0__n264), .A2(ALU_DW_rash_0__n403), .B1(ALU_DW_rash_0__n597), .B2(ALU_DW_rash_0__n492), .Y(
        n659) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U733 ( .A1(ALU_DW_rash_0__n35), .A2(ALU_DW_rash_0__n579), .B1(n1215), .B2(ALU_DW_rash_0__n587), .Y(
        n690) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U734 ( .A1(n969), .A2(ALU_DW_rash_0__n578), .B1(ALU_DW_rash_0__n38), .B2(ALU_DW_rash_0__n587), .Y(
        n691) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U735 ( .A1(n1100), .A2(ALU_DW_rash_0__n577), .B1(ALU_DW_rash_0__n373), .B2(ALU_DW_rash_0__n588), .Y(
        n692) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U736 ( .A1(ALU_DW_rash_0__n507), .A2(ALU_DW_rash_0__n549), .B1(ALU_DW_rash_0__n462), .B2(ALU_DW_rash_0__n408), .C1(
        n479), .C2(ALU_DW_rash_0__n183), .Y(ALU_DW_rash_0__n693) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U737 ( .A1(n1225), .A2(ALU_DW_rash_0__n578), .B1(n1068), .B2(ALU_DW_rash_0__n588), .Y(
        n695) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U738 ( .A1(n969), .A2(ALU_DW_rash_0__n563), .B1(n925), .B2(ALU_DW_rash_0__n553), .Y(
        n696) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U739 ( .A1(ALU_DW_rash_0__n373), .A2(ALU_DW_rash_0__n577), .B1(n1064), .B2(ALU_DW_rash_0__n588), .Y(
        n697) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U740 ( .A1(ALU_DW_rash_0__n454), .A2(ALU_DW_rash_0__n59), .B1(ALU_DW_rash_0__n439), .B2(ALU_DW_rash_0__n489), .Y(ALU_DW_rash_0__n660) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U741 ( .A1(n1215), .A2(ALU_DW_rash_0__n577), .B1(n920), .B2(ALU_DW_rash_0__n588), .Y(
        n698) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U742 ( .A1(ALU_DW_rash_0__n38), .A2(ALU_DW_rash_0__n578), .B1(n1109), .B2(ALU_DW_rash_0__n589), .Y(
        n699) );
  OR3x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U743 ( .A(n798), .B(n888), .C(ALU_DW_rash_0__n278), .Y(ALU_DW_rash_0__n706) );
  OR3x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U744 ( .A(n851), .B(n955), .C(n1056), .Y(ALU_DW_rash_0__n707) );
  OR3x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U745 ( .A(n858), .B(n790), .C(n547), .Y(ALU_DW_rash_0__n708) );
  OR3x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U746 ( .A(n1222), .B(n794), .C(n767), .Y(ALU_DW_rash_0__n709) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U747 ( .A1(ALU_DW_rash_0__n434), .A2(ALU_DW_rash_0__n577), .B1(n973), .B2(ALU_DW_rash_0__n588), .Y(
        n711) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U748 ( .A1(n925), .A2(ALU_DW_rash_0__n72), .B1(n969), .B2(ALU_DW_rash_0__n587), .Y(
        n712) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW_rash_0___U749 ( .A1(ALU_DW_rash_0__n477), .A2(ALU_DW_rash_0__n517), .B1(ALU_DW_rash_0__n509), .B2(ALU_DW_rash_0__n410), .Y(
        n714) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U750 ( .A1(n1160), .A2(ALU_DW_rash_0__n580), .B1(n1100), .B2(ALU_DW_rash_0__n589), .Y(
        n716) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U751 ( .A1(ALU_DW_rash_0__n407), .A2(ALU_DW_rash_0__n580), .B1(n1182), .B2(ALU_DW_rash_0__n589), .Y(
        n717) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U752 ( .A1(ALU_DW_rash_0__n385), .A2(ALU_DW_rash_0__n579), .B1(n1024), .B2(ALU_DW_rash_0__n589), .Y(
        n718) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW_rash_0___U753 ( .A1(ALU_DW_rash_0__n590), .A2(ALU_DW_rash_0__n406), .B1(ALU_DW_rash_0__n578), .B2(n1060), .Y(
        n719) );

 AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U1 ( .A(ID_EX_inst_addr[8]), .B(ALU_DW01_add_0__n99), .Y(ALU_DW01_add_0__n114) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U2 ( .A(ID_EX_inst_addr[26]), .B(ALU_DW01_add_0__n73), .Y(ALU_DW01_add_0__n122) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U3 ( .A(n12), .B(ALU_DW01_add_0__n87), .Y(ALU_DW01_add_0__n140) );
  INVxp33_ASAP7_75t_R ALU___ALU_DW01_add_0___U4 ( .A(n10), .Y(ALU_DW01_add_0__n180) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U5 ( .A(n24), .B(ALU_DW01_add_0__n30), .Y(ALU_DW01_add_0__n124) );
  BUFx4_ASAP7_75t_R ALU___ALU_DW01_add_0___U6 ( .A(ID_EX_inst_addr[0]), .Y(ALU__N323) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_0___U7 ( .A(n25), .Y(ALU_DW01_add_0__n240) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U8 ( .A(n38), .B(n25), .Y(ALU_DW01_add_0__n119) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U9 ( .A(n49), .B(ALU_DW01_add_0__n36), .Y(ALU_DW01_add_0__n123) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U10 ( .A(n21), .B(ALU_DW01_add_0__n118), .Y(ALU_DW01_add_0__n142) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U11 ( .A(n39), .B(ALU_DW01_add_0__n5), .Y(ALU_DW01_add_0__n138) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U12 ( .A(ID_EX_inst_addr[17]), .B(ALU_DW01_add_0__n127), .Y(ALU_DW01_add_0__n145) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U13 ( .A(n69), .B(ALU_DW01_add_0__n110), .Y(ALU_DW01_add_0__n134) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U14 ( .A(ALU_DW01_add_0__ALU_DW01_add_0__n112), .Y(ALU_DW01_add_0__n1) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U15 ( .A(ALU_DW01_add_0__n64), .Y(ALU_DW01_add_0__n2) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U16 ( .A(ALU_DW01_add_0__n64), .Y(ALU_DW01_add_0__n3) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U17 ( .A(ALU_DW01_add_0__n66), .Y(ALU_DW01_add_0__n4) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U18 ( .A(ALU_DW01_add_0__n66), .Y(ALU_DW01_add_0__n5) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U19 ( .A(ALU_DW01_add_0__n120), .Y(ALU_DW01_add_0__n6) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U20 ( .A(ALU_DW01_add_0__n121), .Y(ALU_DW01_add_0__n7) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U21 ( .A(ALU_DW01_add_0__n102), .Y(ALU_DW01_add_0__n8) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U22 ( .A(ALU_DW01_add_0__n137), .Y(ALU_DW01_add_0__n9) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U23 ( .A(ALU_DW01_add_0__n11), .Y(ALU_DW01_add_0__n10) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_0___U24 ( .A(ALU_DW01_add_0__n179), .Y(ALU_DW01_add_0__n11) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U25 ( .A(ALU_DW01_add_0__n182), .Y(ALU_DW01_add_0__n155) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U26 ( .A(ALU_DW01_add_0__n155), .Y(ALU_DW01_add_0__n12) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U27 ( .A(ALU_DW01_add_0__ALU_DW01_add_0__n134), .Y(ALU_DW01_add_0__n13) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U28 ( .A(ALU_DW01_add_0__ALU_DW01_add_0__n146), .Y(ALU_DW01_add_0__n14) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U29 ( .A(ALU_DW01_add_0__n124), .Y(ALU_DW01_add_0__n15) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U30 ( .A(ALU_DW01_add_0__n9), .Y(ALU_DW01_add_0__n16) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U31 ( .A(ALU_DW01_add_0__n16), .Y(ALU_DW01_add_0__n17) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U32 ( .A(ALU_DW01_add_0__n68), .Y(ALU_DW01_add_0__n18) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U33 ( .A(ALU_DW01_add_0__n68), .Y(ALU_DW01_add_0__n19) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U34 ( .A(ALU_DW01_add_0__n147), .Y(ALU_DW01_add_0__n20) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U35 ( .A(ALU_DW01_add_0__n145), .Y(ALU_DW01_add_0__n21) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U36 ( .A(ALU_DW01_add_0__n141), .Y(ALU_DW01_add_0__n22) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_0___U37 ( .A(ALU_DW01_add_0__n139), .Y(ALU_DW01_add_0__n63) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U38 ( .A(ALU_DW01_add_0__n24), .Y(ALU_DW01_add_0__n23) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U39 ( .A(ALU_DW01_add_0__n186), .Y(ALU_DW01_add_0__n24) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_0___U40 ( .A(ALU_DW01_add_0__n23), .Y(ALU_DW01_add_0__n215) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_0___U41 ( .A(ALU_DW01_add_0__n26), .Y(ALU_DW01_add_0__n25) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U42 ( .A(ALU_DW01_add_0__n135), .Y(ALU_DW01_add_0__n26) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U43 ( .A(ALU_DW01_add_0__n105), .Y(ALU_DW01_add_0__n27) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U44 ( .A(ALU_DW01_add_0__n105), .Y(ALU_DW01_add_0__n28) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U45 ( .A(ALU_DW01_add_0__n1), .Y(ALU_DW01_add_0__n29) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U46 ( .A(ALU_DW01_add_0__n29), .Y(ALU_DW01_add_0__n30) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U47 ( .A(ALU_DW01_add_0__n32), .Y(ALU_DW01_add_0__n31) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U48 ( .A(ALU_DW01_add_0__n198), .Y(ALU_DW01_add_0__n32) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_0___U49 ( .A(ALU_DW01_add_0__n34), .Y(ALU_DW01_add_0__n33) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U50 ( .A(ALU_DW01_add_0__n133), .Y(ALU_DW01_add_0__n34) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U51 ( .A(ALU_DW01_add_0__n78), .Y(ALU_DW01_add_0__n35) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U52 ( .A(ALU_DW01_add_0__n78), .Y(ALU_DW01_add_0__n36) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U53 ( .A(ID_EX_inst_addr[11]), .B(ALU_DW01_add_0__n19), .Y(ALU_DW01_add_0__n103) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U54 ( .A(ALU_DW01_add_0__n138), .Y(ALU_DW01_add_0__n37) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U55 ( .A(ALU_DW01_add_0__n37), .Y(ALU_DW01_add_0__n126) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U56 ( .A(ALU_DW01_add_0__n39), .Y(ALU_DW01_add_0__n38) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U57 ( .A(ALU_DW01_add_0__n128), .Y(ALU_DW01_add_0__n39) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U58 ( .A(ALU_DW01_add_0__n42), .Y(ALU_DW01_add_0__n40) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U59 ( .A(ALU_DW01_add_0__n42), .Y(ALU_DW01_add_0__n41) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U60 ( .A(ALU_DW01_add_0__n22), .Y(ALU_DW01_add_0__n42) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U61 ( .A(ALU_DW01_add_0__n15), .Y(ALU_DW01_add_0__n43) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U62 ( .A(ALU_DW01_add_0__n43), .Y(ALU_DW01_add_0__n44) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U63 ( .A(ALU_DW01_add_0__n129), .Y(ALU_DW01_add_0__n45) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U64 ( .A(ALU_DW01_add_0__n119), .Y(ALU_DW01_add_0__n46) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U65 ( .A(ALU_DW01_add_0__n122), .Y(ALU_DW01_add_0__n47) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_0___U66 ( .A(ALU_DW01_add_0__n130), .Y(ALU_DW01_add_0__n77) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U67 ( .A(ALU_DW01_add_0__n49), .Y(ALU_DW01_add_0__n48) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U68 ( .A(ALU_DW01_add_0__n197), .Y(ALU_DW01_add_0__n49) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U69 ( .A(n20), .B(ALU_DW01_add_0__n3), .Y(ALU_DW01_add_0__n113) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U70 ( .A(ALU_DW01_add_0__n52), .Y(ALU_DW01_add_0__n50) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U71 ( .A(ALU_DW01_add_0__n52), .Y(ALU_DW01_add_0__n51) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U72 ( .A(ALU_DW01_add_0__n7), .Y(ALU_DW01_add_0__n52) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U73 ( .A(ALU__n1080), .Y(ALU_DW01_add_0__n53) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U74 ( .A(ALU__n1080), .Y(ALU_DW01_add_0__n54) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U75 ( .A(ALU__n1081), .Y(ALU_DW01_add_0__n55) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U76 ( .A(ALU__n1081), .Y(ALU_DW01_add_0__n56) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U77 ( .A(ALU_DW01_add_0__n157), .Y(ALU__N344) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U78 ( .A(ALU_DW01_add_0__n59), .Y(ALU_DW01_add_0__n58) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U79 ( .A(ALU_DW01_add_0__n194), .Y(ALU_DW01_add_0__n59) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_0___U80 ( .A(ALU_DW01_add_0__n58), .Y(ALU_DW01_add_0__n223) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U81 ( .A(ALU_DW01_add_0__n61), .Y(ALU_DW01_add_0__n60) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U82 ( .A(ALU_DW01_add_0__n195), .Y(ALU_DW01_add_0__n61) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_0___U83 ( .A(ALU_DW01_add_0__n60), .Y(ALU_DW01_add_0__n224) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U84 ( .A(ALU_DW01_add_0__n63), .Y(ALU_DW01_add_0__n62) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U85 ( .A(ALU_DW01_add_0__n62), .Y(ALU_DW01_add_0__n131) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U86 ( .A(ALU_DW01_add_0__n65), .Y(ALU_DW01_add_0__n64) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U87 ( .A(ALU_DW01_add_0__n140), .Y(ALU_DW01_add_0__n65) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U88 ( .A(ALU_DW01_add_0__n67), .Y(ALU_DW01_add_0__n66) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U89 ( .A(ALU_DW01_add_0__n111), .Y(ALU_DW01_add_0__n67) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U90 ( .A(ALU_DW01_add_0__n69), .Y(ALU_DW01_add_0__n68) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U91 ( .A(ALU_DW01_add_0__n142), .Y(ALU_DW01_add_0__n69) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U92 ( .A(ALU_DW01_add_0__n71), .Y(ALU_DW01_add_0__n70) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U93 ( .A(ALU_DW01_add_0__n114), .Y(ALU_DW01_add_0__n71) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U94 ( .A(ALU_DW01_add_0__n8), .Y(ALU_DW01_add_0__n72) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U95 ( .A(ALU_DW01_add_0__n72), .Y(ALU_DW01_add_0__n73) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U96 ( .A(ALU__n1110), .Y(ALU_DW01_add_0__n74) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U97 ( .A(ALU__n1110), .Y(ALU_DW01_add_0__n75) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U98 ( .A(ALU_DW01_add_0__n77), .Y(ALU_DW01_add_0__n76) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U99 ( .A(ALU_DW01_add_0__n76), .Y(ALU_DW01_add_0__n117) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U100 ( .A(ALU_DW01_add_0__n79), .Y(ALU_DW01_add_0__n78) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U101 ( .A(ALU_DW01_add_0__n103), .Y(ALU_DW01_add_0__n79) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U102 ( .A(ALU_DW01_add_0__n82), .Y(ALU_DW01_add_0__n80) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U103 ( .A(ALU_DW01_add_0__n82), .Y(ALU_DW01_add_0__n81) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U104 ( .A(ALU_DW01_add_0__n21), .Y(ALU_DW01_add_0__n82) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U105 ( .A(ALU_DW01_add_0__n85), .Y(ALU_DW01_add_0__n83) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U106 ( .A(ALU_DW01_add_0__n85), .Y(ALU_DW01_add_0__n84) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U107 ( .A(ALU_DW01_add_0__n14), .Y(ALU_DW01_add_0__n85) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U108 ( .A(ALU_DW01_add_0__n88), .Y(ALU_DW01_add_0__n86) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U109 ( .A(ALU_DW01_add_0__n88), .Y(ALU_DW01_add_0__n87) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U110 ( .A(ALU_DW01_add_0__n47), .Y(ALU_DW01_add_0__n88) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U111 ( .A(ALU_DW01_add_0__n13), .Y(ALU_DW01_add_0__n89) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U112 ( .A(ALU_DW01_add_0__n89), .Y(ALU_DW01_add_0__n90) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U113 ( .A(n2), .B(ALU_DW01_add_0__n90), .Y(ALU_DW01_add_0__n141) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U114 ( .A(ALU_DW01_add_0__n92), .Y(ALU_DW01_add_0__n91) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U115 ( .A(ALU_DW01_add_0__n46), .Y(ALU_DW01_add_0__n92) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U116 ( .A(n27), .B(ALU_DW01_add_0__n92), .Y(ALU_DW01_add_0__n137) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U117 ( .A(ALU_DW01_add_0__n94), .Y(ALU_DW01_add_0__n93) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U118 ( .A(ALU_DW01_add_0__n113), .Y(ALU_DW01_add_0__n94) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U119 ( .A(ALU_DW01_add_0__n97), .Y(ALU_DW01_add_0__n95) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U120 ( .A(ALU_DW01_add_0__n97), .Y(ALU_DW01_add_0__n96) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U121 ( .A(ALU_DW01_add_0__n6), .Y(ALU_DW01_add_0__n97) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U122 ( .A(ALU_DW01_add_0__n20), .Y(ALU_DW01_add_0__n98) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U123 ( .A(ALU_DW01_add_0__n98), .Y(ALU_DW01_add_0__n99) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U124 ( .A(ALU_DW01_add_0__n54), .B(ALU_DW01_add_0__n44), .Y(ALU_DW01_add_0__n147) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U125 ( .A(ALU__n1166), .Y(ALU_DW01_add_0__n100) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U126 ( .A(ALU__n1166), .Y(ALU_DW01_add_0__n101) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U127 ( .A(n1), .B(ALU_DW01_add_0__n28), .Y(ALU_DW01_add_0__n102) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U128 ( .A(ALU_DW01_add_0__n240), .Y(ALU__N325) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U129 ( .A(ALU_DW01_add_0__n106), .Y(ALU_DW01_add_0__n105) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U130 ( .A(ALU_DW01_add_0__n25), .Y(ALU_DW01_add_0__n106) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U131 ( .A(inst_addr[23]), .B(ALU_DW01_add_0__n51), .Y(ALU_DW01_add_0__n128) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U132 ( .A(ALU_DW01_add_0__n108), .Y(ALU_DW01_add_0__n107) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U133 ( .A(ALU_DW01_add_0__n123), .Y(ALU_DW01_add_0__n108) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U134 ( .A(ALU_DW01_add_0__n45), .Y(ALU_DW01_add_0__n109) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U135 ( .A(ALU_DW01_add_0__n109), .Y(ALU_DW01_add_0__n110) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U136 ( .A(ID_EX_inst_addr[19]), .B(ALU_DW01_add_0__n96), .Y(ALU_DW01_add_0__n129) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U137 ( .A(ALU__n1318), .B(ALU_DW01_add_0__n84), .Y(ALU_DW01_add_0__n111) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U138 ( .A(ALU_DW01_add_0__n56), .B(ALU_DW01_add_0__n17), .Y(ALU_DW01_add_0__n112) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_0___U139 ( .A(ALU_DW01_add_0__n116), .Y(ALU_DW01_add_0__n115) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U140 ( .A(ALU_DW01_add_0__n33), .Y(ALU_DW01_add_0__n116) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U141 ( .A(ALU_DW01_add_0__n117), .Y(ALU_DW01_add_0__n118) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U142 ( .A(n4), .B(ALU_DW01_add_0__n81), .Y(ALU_DW01_add_0__n120) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U143 ( .A(ALU_DW01_add_0__n75), .B(ALU_DW01_add_0__n41), .Y(ALU_DW01_add_0__n121) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U144 ( .A(ALU_DW01_add_0__n183), .Y(ALU_DW01_add_0__n125) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_0___U145 ( .A(ALU_DW01_add_0__n125), .Y(ALU_DW01_add_0__n212) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U146 ( .A(ALU_DW01_add_0__n126), .Y(ALU_DW01_add_0__n127) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U147 ( .A(n15), .B(ALU_DW01_add_0__n70), .Y(ALU_DW01_add_0__n130) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_0___U148 ( .A(ALU_DW01_add_0__n151), .Y(ALU_DW01_add_0__n150) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_0___U149 ( .A(ALU_DW01_add_0__n131), .Y(ALU_DW01_add_0__n132) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_0___U150 ( .A(ALU_DW01_add_0__n101), .B(ALU_DW01_add_0__n132), .Y(ALU_DW01_add_0__n146) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U151 ( .A(inst_addr[29]), .B(ALU_DW01_add_0__n93), .Y(ALU_DW01_add_0__n133) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U152 ( .A(inst_addr[24]), .B(ALU_DW01_add_0__n38), .Y(ALU_DW01_add_0__n135) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U153 ( .A(ALU_DW01_add_0__n210), .Y(ALU_DW01_add_0__n239) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U154 ( .A(ALU_DW01_add_0__n239), .Y(ALU__N326) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U155 ( .A(n17), .B(ALU_DW01_add_0__n107), .Y(ALU_DW01_add_0__n139) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U156 ( .A(ALU_DW01_add_0__n188), .Y(ALU_DW01_add_0__n217) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U157 ( .A(ALU_DW01_add_0__n217), .Y(ALU__N348) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U158 ( .A(ALU_DW01_add_0__n193), .Y(ALU_DW01_add_0__n222) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U159 ( .A(ALU_DW01_add_0__n222), .Y(ALU__N343) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_0___U160 ( .A(ALU_DW01_add_0__n180), .Y(ALU__N324) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U161 ( .A(ALU_DW01_add_0__n212), .Y(ALU__N353) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U162 ( .A(ALU_DW01_add_0__n214), .Y(ALU__N351) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U163 ( .A(ALU_DW01_add_0__n185), .Y(ALU_DW01_add_0__n151) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_0___U164 ( .A(ALU_DW01_add_0__n150), .Y(ALU_DW01_add_0__n214) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U165 ( .A(ALU_DW01_add_0__n184), .Y(ALU_DW01_add_0__n213) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U166 ( .A(ALU_DW01_add_0__n213), .Y(ALU__N352) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U167 ( .A(ALU_DW01_add_0__n181), .Y(ALU_DW01_add_0__n211) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U168 ( .A(ALU_DW01_add_0__n211), .Y(ALU__N354) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U169 ( .A(ALU_DW01_add_0__n12), .Y(ALU_DW01_add_0__n179) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U170 ( .A(ALU_DW01_add_0__n10), .Y(ALU_DW01_add_0__n154) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U171 ( .A(inst_addr[30]), .B(ALU_DW01_add_0__n115), .Y(ALU_DW01_add_0__n182) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U172 ( .A(inst_addr[31]), .B(ALU_DW01_add_0__n154), .Y(ALU_DW01_add_0__n181) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U173 ( .A(ALU_DW01_add_0__n187), .Y(ALU_DW01_add_0__n216) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U174 ( .A(ALU_DW01_add_0__n216), .Y(ALU__N349) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U175 ( .A(ALU_DW01_add_0__n72), .B(ID_EX_inst_addr[26]), .Y(ALU_DW01_add_0__n187) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U176 ( .A(ALU_DW01_add_0__n192), .Y(ALU_DW01_add_0__n221) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U177 ( .A(ALU_DW01_add_0__n221), .Y(ALU_DW01_add_0__n157) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U178 ( .A(ALU_DW01_add_0__n89), .B(n2), .Y(ALU_DW01_add_0__n192) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U179 ( .A(ALU_DW01_add_0__n201), .Y(ALU_DW01_add_0__n230) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U180 ( .A(ALU_DW01_add_0__n230), .Y(ALU__N335) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U181 ( .A(ALU_DW01_add_0__n35), .B(n49), .Y(ALU_DW01_add_0__n201) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U182 ( .A(ALU_DW01_add_0__n209), .Y(ALU_DW01_add_0__n238) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U183 ( .A(ALU_DW01_add_0__n238), .Y(ALU__N327) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U184 ( .A(ALU_DW01_add_0__n91), .B(n27), .Y(ALU_DW01_add_0__n209) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U185 ( .A(ALU_DW01_add_0__n215), .Y(ALU__N350) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U186 ( .A(ALU_DW01_add_0__n86), .B(n12), .Y(ALU_DW01_add_0__n186) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U187 ( .A(ALU_DW01_add_0__n189), .Y(ALU_DW01_add_0__n218) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U188 ( .A(ALU_DW01_add_0__n218), .Y(ALU__N347) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U189 ( .A(ALU_DW01_add_0__n38), .B(inst_addr[24]), .Y(ALU_DW01_add_0__n189) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U190 ( .A(ALU_DW01_add_0__n190), .Y(ALU_DW01_add_0__n219) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U191 ( .A(ALU_DW01_add_0__n219), .Y(ALU__N346) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U192 ( .A(ALU_DW01_add_0__n50), .B(inst_addr[23]), .Y(ALU_DW01_add_0__n190) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U193 ( .A(ALU_DW01_add_0__n191), .Y(ALU_DW01_add_0__n220) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U194 ( .A(ALU_DW01_add_0__n220), .Y(ALU__N345) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U195 ( .A(ALU_DW01_add_0__n40), .B(ALU_DW01_add_0__n74), .Y(ALU_DW01_add_0__n191) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U196 ( .A(ALU_DW01_add_0__n223), .Y(ALU__N342) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U197 ( .A(ALU_DW01_add_0__n95), .B(ID_EX_inst_addr[19]), .Y(ALU_DW01_add_0__n194) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U198 ( .A(ALU_DW01_add_0__n224), .Y(ALU__N341) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U199 ( .A(ALU_DW01_add_0__n80), .B(n4), .Y(ALU_DW01_add_0__n195) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U200 ( .A(ALU_DW01_add_0__n196), .Y(ALU_DW01_add_0__n225) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U201 ( .A(ALU_DW01_add_0__n225), .Y(ALU__N340) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U202 ( .A(ALU_DW01_add_0__n126), .B(ID_EX_inst_addr[17]), .Y(ALU_DW01_add_0__n196) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U203 ( .A(ALU_DW01_add_0__n48), .Y(ALU_DW01_add_0__n226) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U204 ( .A(ALU_DW01_add_0__n226), .Y(ALU__N339) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U205 ( .A(ALU_DW01_add_0__n4), .B(n39), .Y(ALU_DW01_add_0__n197) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U206 ( .A(ALU_DW01_add_0__n31), .Y(ALU_DW01_add_0__n227) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U207 ( .A(ALU_DW01_add_0__n227), .Y(ALU__N338) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U208 ( .A(ALU_DW01_add_0__n83), .B(ALU__n1318), .Y(ALU_DW01_add_0__n198) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U209 ( .A(ALU_DW01_add_0__n199), .Y(ALU_DW01_add_0__n228) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U210 ( .A(ALU_DW01_add_0__n228), .Y(ALU__N337) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U211 ( .A(ALU_DW01_add_0__n131), .B(ALU_DW01_add_0__n100), .Y(ALU_DW01_add_0__n199) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U212 ( .A(ALU_DW01_add_0__n200), .Y(ALU_DW01_add_0__n229) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U213 ( .A(ALU_DW01_add_0__n229), .Y(ALU__N336) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U214 ( .A(ALU_DW01_add_0__n107), .B(n17), .Y(ALU_DW01_add_0__n200) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U215 ( .A(ALU_DW01_add_0__n202), .Y(ALU_DW01_add_0__n231) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U216 ( .A(ALU_DW01_add_0__n231), .Y(ALU__N334) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U217 ( .A(ALU_DW01_add_0__n18), .B(ID_EX_inst_addr[11]), .Y(ALU_DW01_add_0__n202) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U218 ( .A(ALU_DW01_add_0__n203), .Y(ALU_DW01_add_0__n232) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U219 ( .A(ALU_DW01_add_0__n232), .Y(ALU__N333) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U220 ( .A(ALU_DW01_add_0__n117), .B(n21), .Y(ALU_DW01_add_0__n203) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U221 ( .A(ALU_DW01_add_0__n204), .Y(ALU_DW01_add_0__n233) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U222 ( .A(ALU_DW01_add_0__n233), .Y(ALU__N332) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U223 ( .A(ALU_DW01_add_0__n70), .B(n15), .Y(ALU_DW01_add_0__n204) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U224 ( .A(ALU_DW01_add_0__n205), .Y(ALU_DW01_add_0__n234) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U225 ( .A(ALU_DW01_add_0__n234), .Y(ALU__N331) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U226 ( .A(ALU_DW01_add_0__n98), .B(ID_EX_inst_addr[8]), .Y(ALU_DW01_add_0__n205) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U227 ( .A(ALU_DW01_add_0__n206), .Y(ALU_DW01_add_0__n235) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U228 ( .A(ALU_DW01_add_0__n235), .Y(ALU__N330) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U229 ( .A(ALU_DW01_add_0__n43), .B(ALU_DW01_add_0__n53), .Y(ALU_DW01_add_0__n206) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U230 ( .A(ALU_DW01_add_0__n207), .Y(ALU_DW01_add_0__n236) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U231 ( .A(ALU_DW01_add_0__n236), .Y(ALU__N329) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U232 ( .A(ALU_DW01_add_0__n29), .B(n24), .Y(ALU_DW01_add_0__n207) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_0___U233 ( .A(ALU_DW01_add_0__n208), .Y(ALU_DW01_add_0__n237) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_0___U234 ( .A(ALU_DW01_add_0__n237), .Y(ALU__N328) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U235 ( .A(ALU_DW01_add_0__n16), .B(ALU_DW01_add_0__n55), .Y(ALU_DW01_add_0__n208) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U236 ( .A(ALU_DW01_add_0__n27), .B(n1), .Y(ALU_DW01_add_0__n188) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U237 ( .A(ALU_DW01_add_0__n109), .B(n69), .Y(ALU_DW01_add_0__n193) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U238 ( .A(ALU_DW01_add_0__n93), .B(inst_addr[29]), .Y(ALU_DW01_add_0__n184) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U239 ( .A(ALU_DW01_add_0__n2), .B(n20), .Y(ALU_DW01_add_0__n185) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U240 ( .A(ALU_DW01_add_0__n115), .B(inst_addr[30]), .Y(ALU_DW01_add_0__n183) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_0___U241 ( .A(n25), .B(n38), .Y(ALU_DW01_add_0__n210) );

  INVxp33_ASAP7_75t_R ALU___ALU_DW01_ash_0___U3 ( .A(ALU_DW01_ash_0__n1), .Y(ALU_DW01_ash_0__n818) );
  NOR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U4 ( .A(ALU_DW01_ash_0__n601), .B(ALU_DW01_ash_0__n3), .Y(ALU_DW01_ash_0__n2) );
  NOR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U5 ( .A(ALU_DW01_ash_0__n609), .B(ALU_DW01_ash_0__n197), .Y(ALU_DW01_ash_0__n4) );
  NOR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U6 ( .A(ALU_DW01_ash_0__n131), .B(ALU_DW01_ash_0__ALU_DW01_ash_0__n539), .Y(ALU_DW01_ash_0__n5) );
  NOR2xp67_ASAP7_75t_R ALU___ALU_DW01_ash_0___U7 ( .A(ALU_DW01_ash_0__n5), .B(ALU_DW01_ash_0__n6), .Y(ALU_DW01_ash_0__n1) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_ash_0___U8 ( .A(ALU_DW01_ash_0__n463), .B(ALU__n901), .Y(ALU_DW01_ash_0__n7) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U9 ( .A(ALU_DW01_ash_0__n7), .Y(ALU_DW01_ash_0__n3) );
  NOR2x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U10 ( .A(ALU_DW01_ash_0__n2), .B(ALU_DW01_ash_0__n4), .Y(ALU_DW01_ash_0__n8) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U11 ( .A(ALU_DW01_ash_0__n8), .Y(ALU_DW01_ash_0__n6) );
  CKINVDCx6p67_ASAP7_75t_R ALU___ALU_DW01_ash_0___U12 ( .A(ALU_DW01_ash_0__n266), .Y(ALU_DW01_ash_0__n609) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U13 ( .A(ALU_DW01_ash_0__n393), .Y(ALU_DW01_ash_0__n9) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U14 ( .A(ALU_DW01_ash_0__n651), .Y(ALU_DW01_ash_0__n10) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U15 ( .A(ALU_DW01_ash_0__n654), .Y(ALU_DW01_ash_0__n11) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U16 ( .A(ALU_DW01_ash_0__n13), .Y(ALU_DW01_ash_0__n12) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U17 ( .A(ALU_DW01_ash_0__n299), .Y(ALU_DW01_ash_0__n13) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U18 ( .A(ALU_DW01_ash_0__n34), .Y(ALU_DW01_ash_0__n528) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U19 ( .A(ALU_DW01_ash_0__n300), .Y(ALU_DW01_ash_0__n299) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U20 ( .A(ALU_DW01_ash_0__n433), .Y(ALU_DW01_ash_0__n14) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U21 ( .A(ALU_DW01_ash_0__n644), .Y(ALU_DW01_ash_0__n15) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U22 ( .A(ALU_DW01_ash_0__n743), .Y(ALU_DW01_ash_0__n16) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U23 ( .A(ALU_DW01_ash_0__n656), .Y(ALU_DW01_ash_0__n17) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U24 ( .A(ALU_DW01_ash_0__n404), .Y(ALU_DW01_ash_0__n18) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U25 ( .A(ALU_DW01_ash_0__n20), .Y(ALU_DW01_ash_0__n19) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U26 ( .A(ALU_DW01_ash_0__n11), .Y(ALU_DW01_ash_0__n20) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U27 ( .A(ALU_DW01_ash_0__n19), .Y(ALU_DW01_ash_0__n405) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U28 ( .A(ALU_DW01_ash_0__n405), .Y(ALU_DW01_ash_0__n21) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U29 ( .A(ALU_DW01_ash_0__n657), .Y(ALU_DW01_ash_0__n22) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U30 ( .A(ALU_DW01_ash_0__n658), .Y(ALU_DW01_ash_0__n23) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U31 ( .A(ALU_DW01_ash_0__n659), .Y(ALU_DW01_ash_0__n24) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U32 ( .A(ALU_DW01_ash_0__n288), .Y(ALU_DW01_ash_0__n33) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U33 ( .A(ALU__n73), .Y(ALU_DW01_ash_0__n25) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U34 ( .A(ALU_DW01_ash_0__n673), .Y(ALU_DW01_ash_0__n26) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U35 ( .A(ALU_DW01_ash_0__n673), .Y(ALU_DW01_ash_0__n27) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U36 ( .A(ALU_DW01_ash_0__n676), .Y(ALU_DW01_ash_0__n28) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U37 ( .A(ALU_DW01_ash_0__n676), .Y(ALU_DW01_ash_0__n29) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U38 ( .A(ALU__n80), .Y(ALU_DW01_ash_0__n30) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U39 ( .A(ALU_DW01_ash_0__n32), .Y(ALU_DW01_ash_0__n31) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U40 ( .A(ALU_DW01_ash_0__n865), .Y(ALU_DW01_ash_0__n32) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U41 ( .A(ALU_DW01_ash_0__n31), .Y(ALU_DW01_ash_0__n77) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U42 ( .A(ALU_DW01_ash_0__n36), .Y(ALU_DW01_ash_0__n34) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U43 ( .A(ALU_DW01_ash_0__n37), .Y(ALU_DW01_ash_0__n35) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U44 ( .A(ALU_DW01_ash_0__ALU_DW01_ash_0__n368), .Y(ALU_DW01_ash_0__n36) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U45 ( .A(ALU_DW01_ash_0__n368), .Y(ALU_DW01_ash_0__n37) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U46 ( .A(ALU_DW01_ash_0__n857), .Y(ALU_DW01_ash_0__n38) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U47 ( .A(ALU_DW01_ash_0__n38), .Y(ALU_DW01_ash_0__n41) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U48 ( .A(ALU_DW01_ash_0__n691), .Y(ALU_DW01_ash_0__n39) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U49 ( .A(ALU_DW01_ash_0__n691), .Y(ALU_DW01_ash_0__n40) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U50 ( .A(ALU_DW01_ash_0__n531), .Y(ALU_DW01_ash_0__n691) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U51 ( .A(ALU_DW01_ash_0__n728), .Y(ALU_DW01_ash_0__n42) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U52 ( .A(ALU_DW01_ash_0__n728), .Y(ALU_DW01_ash_0__n43) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U53 ( .A(ALU_DW01_ash_0__n674), .Y(ALU_DW01_ash_0__n44) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U54 ( .A(ALU_DW01_ash_0__n674), .Y(ALU_DW01_ash_0__n45) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U55 ( .A(ALU_DW01_ash_0__n50), .Y(ALU_DW01_ash_0__n46) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U56 ( .A(ALU_DW01_ash_0__n693), .Y(ALU_DW01_ash_0__n686) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U57 ( .A(ALU_DW01_ash_0__n287), .Y(ALU_DW01_ash_0__n693) );
  INVx5_ASAP7_75t_R ALU___ALU_DW01_ash_0___U58 ( .A(ALU_DW01_ash_0__n532), .Y(ALU_DW01_ash_0__n688) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U59 ( .A(ALU_DW01_ash_0__n615), .Y(ALU_DW01_ash_0__n685) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U60 ( .A(n1020), .Y(ALU_DW01_ash_0__n47) );
  AO22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U61 ( .A1(ALU_DW01_ash_0__n140), .A2(ALU_DW01_ash_0__n721), .B1(n1020), .B2(ALU_DW01_ash_0__n701), .Y(
        n832) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U62 ( .A(ALU_DW01_ash_0__n858), .Y(ALU_DW01_ash_0__n48) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U63 ( .A(ALU_DW01_ash_0__n53), .Y(ALU_DW01_ash_0__n49) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U64 ( .A(ALU_DW01_ash_0__n59), .Y(ALU_DW01_ash_0__n50) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U65 ( .A(ALU_DW01_ash_0__n349), .Y(ALU_DW01_ash_0__n51) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U66 ( .A(ALU_DW01_ash_0__n860), .Y(ALU_DW01_ash_0__n52) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U67 ( .A(ALU_DW01_ash_0__n64), .Y(ALU_DW01_ash_0__n53) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U68 ( .A(ALU_DW01_ash_0__n130), .Y(ALU_DW01_ash_0__n54) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U69 ( .A(ALU_DW01_ash_0__n112), .Y(ALU_DW01_ash_0__n55) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U70 ( .A(ALU_DW01_ash_0__n863), .Y(ALU_DW01_ash_0__n56) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U71 ( .A(ALU_DW01_ash_0__n56), .Y(ALU_DW01_ash_0__n70) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U72 ( .A(ALU_DW01_ash_0__n58), .Y(ALU_DW01_ash_0__n57) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U73 ( .A(ALU_DW01_ash_0__n861), .Y(ALU_DW01_ash_0__n58) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U74 ( .A(ALU_DW01_ash_0__n72), .Y(ALU_DW01_ash_0__n59) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U75 ( .A(ALU_DW01_ash_0__n623), .Y(ALU_DW01_ash_0__n60) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U76 ( .A(ALU_DW01_ash_0__n62), .Y(ALU_DW01_ash_0__n61) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U77 ( .A(ALU_DW01_ash_0__n859), .Y(ALU_DW01_ash_0__n62) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U78 ( .A(ALU_DW01_ash_0__n862), .Y(ALU_DW01_ash_0__n63) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U79 ( .A(ALU_DW01_ash_0__n78), .Y(ALU_DW01_ash_0__n64) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U80 ( .A(ALU_DW01_ash_0__n49), .Y(ALU_DW01_ash_0__n65) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U81 ( .A(ALU_DW01_ash_0__n377), .Y(ALU_DW01_ash_0__n66) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U82 ( .A(ALU_DW01_ash_0__n778), .Y(ALU_DW01_ash_0__n67) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U83 ( .A(ALU_DW01_ash_0__n260), .Y(ALU_DW01_ash_0__n68) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U84 ( .A(ALU_DW01_ash_0__n75), .Y(ALU_DW01_ash_0__n69) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U85 ( .A(ALU_DW01_ash_0__n736), .Y(ALU_DW01_ash_0__n71) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U86 ( .A(ALU_DW01_ash_0__n209), .Y(ALU_DW01_ash_0__n72) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U87 ( .A(ALU_DW01_ash_0__n81), .Y(ALU_DW01_ash_0__n73) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U88 ( .A(ALU_DW01_ash_0__n587), .Y(ALU_DW01_ash_0__n631) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U89 ( .A(ALU_DW01_ash_0__n104), .Y(ALU_DW01_ash_0__n74) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U90 ( .A(ALU_DW01_ash_0__n738), .Y(ALU_DW01_ash_0__n75) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U91 ( .A(ALU_DW01_ash_0__n576), .Y(ALU_DW01_ash_0__n575) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U92 ( .A(ALU_DW01_ash_0__n69), .Y(ALU_DW01_ash_0__n576) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U93 ( .A(ALU__n368), .Y(ALU_DW01_ash_0__n76) );
  CKINVDCx16_ASAP7_75t_R ALU___ALU_DW01_ash_0___U94 ( .A(ALU_DW01_ash_0__n689), .Y(ALU_DW01_ash_0__n687) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U95 ( .A(ALU_DW01_ash_0__n729), .Y(ALU_DW01_ash_0__n78) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U96 ( .A(ALU_DW01_ash_0__n851), .Y(ALU_DW01_ash_0__n79) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U97 ( .A(ALU_DW01_ash_0__n91), .Y(ALU_DW01_ash_0__n80) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U98 ( .A(ALU_DW01_ash_0__n739), .Y(ALU_DW01_ash_0__n81) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U99 ( .A(ALU_DW01_ash_0__n356), .Y(ALU_DW01_ash_0__n565) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U100 ( .A(ALU_DW01_ash_0__n600), .Y(ALU_DW01_ash_0__n599) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U101 ( .A(ALU_DW01_ash_0__n73), .Y(ALU_DW01_ash_0__n600) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U102 ( .A(ALU_DW01_ash_0__n830), .Y(ALU_DW01_ash_0__n82) );
  CKINVDCx8_ASAP7_75t_R ALU___ALU_DW01_ash_0___U103 ( .A(ALU_DW01_ash_0__n181), .Y(ALU_DW01_ash_0__n551) );
  CKINVDCx8_ASAP7_75t_R ALU___ALU_DW01_ash_0___U104 ( .A(ALU_DW01_ash_0__n166), .Y(ALU_DW01_ash_0__n607) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U105 ( .A(ALU_DW01_ash_0__n167), .Y(ALU_DW01_ash_0__n166) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U106 ( .A(ALU_DW01_ash_0__n745), .Y(ALU_DW01_ash_0__n83) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U107 ( .A(ALU_DW01_ash_0__n805), .Y(ALU_DW01_ash_0__n84) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U108 ( .A(ALU_DW01_ash_0__n86), .Y(ALU_DW01_ash_0__n85) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U109 ( .A(ALU_DW01_ash_0__n781), .Y(ALU_DW01_ash_0__n86) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U110 ( .A(ALU_DW01_ash_0__n866), .Y(ALU_DW01_ash_0__n87) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U111 ( .A(ALU_DW01_ash_0__n89), .Y(ALU_DW01_ash_0__n88) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U112 ( .A(ALU_DW01_ash_0__n774), .Y(ALU_DW01_ash_0__n89) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U113 ( .A1(ALU_DW01_ash_0__n667), .A2(n1068), .B1(ALU_DW01_ash_0__n680), .B2(ALU_DW01_ash_0__n190), .C(
        n510), .Y(ALU_DW01_ash_0__n774) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U114 ( .A(ALU_DW01_ash_0__n235), .Y(ALU__N271) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U115 ( .A(ALU_DW01_ash_0__n740), .Y(ALU_DW01_ash_0__n91) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U116 ( .A(ALU_DW01_ash_0__n389), .Y(ALU_DW01_ash_0__n388) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U117 ( .A(ALU_DW01_ash_0__n80), .Y(ALU_DW01_ash_0__n389) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U118 ( .A(ALU_DW01_ash_0__n494), .Y(ALU_DW01_ash_0__n340) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U119 ( .A(ALU_DW01_ash_0__n239), .Y(ALU_DW01_ash_0__n92) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U120 ( .A(ALU_DW01_ash_0__n94), .Y(ALU_DW01_ash_0__n93) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U121 ( .A(ALU_DW01_ash_0__n755), .Y(ALU_DW01_ash_0__n94) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U122 ( .A1(ALU_DW01_ash_0__n660), .A2(n1100), .B1(ALU_DW01_ash_0__n679), .B2(n1160), .C(
        n505), .Y(ALU_DW01_ash_0__n755) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U123 ( .A(ALU_DW01_ash_0__n93), .Y(ALU_DW01_ash_0__n165) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U124 ( .A(ALU_DW01_ash_0__n129), .Y(ALU_DW01_ash_0__n95) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U125 ( .A(ALU_DW01_ash_0__n776), .Y(ALU_DW01_ash_0__n96) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U126 ( .A1(ALU_DW01_ash_0__n661), .A2(n1064), .B1(ALU_DW01_ash_0__n680), .B2(ALU_DW01_ash_0__n486), .C(
        n424), .Y(ALU_DW01_ash_0__n776) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U127 ( .A(ALU_DW01_ash_0__n864), .Y(ALU_DW01_ash_0__n97) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U128 ( .A(ALU_DW01_ash_0__n99), .Y(ALU_DW01_ash_0__n98) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U129 ( .A(ALU_DW01_ash_0__n867), .Y(ALU_DW01_ash_0__n99) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U130 ( .A(ALU_DW01_ash_0__n101), .Y(ALU_DW01_ash_0__n100) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U131 ( .A(ALU_DW01_ash_0__n804), .Y(ALU_DW01_ash_0__n101) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U132 ( .A1(ALU_DW01_ash_0__n667), .A2(n1060), .B1(ALU_DW01_ash_0__n684), .B2(ALU_DW01_ash_0__n457), .C(
        n523), .Y(ALU_DW01_ash_0__n804) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U133 ( .A(ALU__n336), .Y(ALU_DW01_ash_0__n102) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U134 ( .A(ALU_DW01_ash_0__n272), .Y(ALU_DW01_ash_0__n103) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U135 ( .A(ALU_DW01_ash_0__n737), .Y(ALU_DW01_ash_0__n104) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U136 ( .A(ALU_DW01_ash_0__n482), .Y(ALU_DW01_ash_0__n481) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U137 ( .A(ALU_DW01_ash_0__n74), .Y(ALU_DW01_ash_0__n482) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U138 ( .A(ALU_DW01_ash_0__n106), .Y(ALU_DW01_ash_0__n105) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U139 ( .A(ALU_DW01_ash_0__n83), .Y(ALU_DW01_ash_0__n106) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U140 ( .A1(ALU_DW01_ash_0__n454), .A2(ALU_DW01_ash_0__n663), .B1(ALU_DW01_ash_0__n392), .B2(ALU_DW01_ash_0__n687), .C(
        n499), .Y(ALU_DW01_ash_0__n745) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U141 ( .A(ALU_DW01_ash_0__n773), .Y(ALU_DW01_ash_0__n107) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U142 ( .A(ALU_DW01_ash_0__n109), .Y(ALU_DW01_ash_0__n108) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U143 ( .A(ALU_DW01_ash_0__n771), .Y(ALU_DW01_ash_0__n109) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U144 ( .A(ALU_DW01_ash_0__n111), .Y(ALU_DW01_ash_0__n110) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U145 ( .A(ALU_DW01_ash_0__n751), .Y(ALU_DW01_ash_0__n111) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U146 ( .A1(ALU_DW01_ash_0__n662), .A2(n1024), .B1(ALU_DW01_ash_0__n680), .B2(ALU_DW01_ash_0__n502), .C(
        n475), .Y(ALU_DW01_ash_0__n751) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U147 ( .A(ALU_DW01_ash_0__n113), .Y(ALU_DW01_ash_0__n112) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U148 ( .A(ALU_DW01_ash_0__n100), .Y(ALU_DW01_ash_0__n113) );
  AO22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U149 ( .A1(ALU_DW01_ash_0__n726), .A2(n1015), .B1(ALU_DW01_ash_0__n705), .B2(ALU_DW01_ash_0__n533), .Y(
        n839) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U150 ( .A(ALU_DW01_ash_0__n55), .Y(ALU_DW01_ash_0__n522) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U151 ( .A(ALU_DW01_ash_0__n116), .Y(ALU_DW01_ash_0__n114) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U152 ( .A(ALU_DW01_ash_0__n116), .Y(ALU_DW01_ash_0__n115) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U153 ( .A(ALU_DW01_ash_0__n14), .Y(ALU_DW01_ash_0__n116) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U154 ( .A(ALU_DW01_ash_0__n640), .Y(ALU_DW01_ash_0__n117) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U155 ( .A(ALU_DW01_ash_0__n641), .Y(ALU_DW01_ash_0__n118) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U156 ( .A(ALU_DW01_ash_0__n120), .Y(ALU_DW01_ash_0__n119) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U157 ( .A(ALU_DW01_ash_0__n642), .Y(ALU_DW01_ash_0__n120) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U158 ( .A(ALU_DW01_ash_0__n122), .Y(ALU_DW01_ash_0__n121) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U159 ( .A(ALU_DW01_ash_0__n15), .Y(ALU_DW01_ash_0__n122) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U160 ( .A(ALU_DW01_ash_0__n121), .Y(ALU_DW01_ash_0__n437) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U161 ( .A(ALU_DW01_ash_0__n437), .Y(ALU_DW01_ash_0__n123) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U162 ( .A(ALU_DW01_ash_0__n834), .Y(ALU_DW01_ash_0__n438) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U163 ( .A(ALU_DW01_ash_0__n438), .Y(ALU_DW01_ash_0__n124) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U164 ( .A(ALU_DW01_ash_0__n645), .Y(ALU_DW01_ash_0__n125) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U165 ( .A(ALU_DW01_ash_0__n436), .B(ALU_DW01_ash_0__n643), .Y(ALU_DW01_ash_0__n433) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U166 ( .A(ALU_DW01_ash_0__n710), .Y(ALU_DW01_ash_0__n702) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U167 ( .A(ALU_DW01_ash_0__n850), .Y(ALU_DW01_ash_0__n126) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U168 ( .A(ALU_DW01_ash_0__n607), .Y(ALU_DW01_ash_0__n732) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U169 ( .A(ALU_DW01_ash_0__n300), .Y(ALU_DW01_ash_0__n301) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U170 ( .A(ALU_DW01_ash_0__n749), .Y(ALU_DW01_ash_0__n127) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U171 ( .A(ALU_DW01_ash_0__n95), .Y(ALU_DW01_ash_0__n128) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U172 ( .A(ALU_DW01_ash_0__n96), .Y(ALU_DW01_ash_0__n129) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U173 ( .A(ALU_DW01_ash_0__n128), .Y(ALU_DW01_ash_0__n426) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U174 ( .A(ALU_DW01_ash_0__n134), .Y(ALU_DW01_ash_0__n355) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U175 ( .A(ALU_DW01_ash_0__n355), .Y(ALU_DW01_ash_0__n130) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U176 ( .A(ALU_DW01_ash_0__n352), .Y(ALU_DW01_ash_0__n131) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U177 ( .A(ALU_DW01_ash_0__n633), .Y(ALU_DW01_ash_0__n132) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U178 ( .A(ALU_DW01_ash_0__n634), .Y(ALU_DW01_ash_0__n133) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U179 ( .A(ALU_DW01_ash_0__n135), .Y(ALU_DW01_ash_0__n134) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U180 ( .A(ALU_DW01_ash_0__n637), .Y(ALU_DW01_ash_0__n135) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U181 ( .A(ALU_DW01_ash_0__n158), .Y(ALU_DW01_ash_0__n136) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U182 ( .A(ALU_DW01_ash_0__n764), .Y(ALU_DW01_ash_0__n137) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U183 ( .A(ALU_DW01_ash_0__n139), .Y(ALU_DW01_ash_0__n138) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U184 ( .A(ALU_DW01_ash_0__n762), .Y(ALU_DW01_ash_0__n139) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U185 ( .A(n1109), .Y(ALU_DW01_ash_0__n140) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U186 ( .A(n1109), .Y(ALU_DW01_ash_0__n141) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U187 ( .A(n1109), .Y(ALU_DW01_ash_0__n142) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U188 ( .A(n1109), .Y(ALU_DW01_ash_0__n143) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U189 ( .A(ALU_DW01_ash_0__n146), .Y(ALU_DW01_ash_0__n144) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U190 ( .A(ALU_DW01_ash_0__n146), .Y(ALU_DW01_ash_0__n145) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U191 ( .A(ALU_DW01_ash_0__n9), .Y(ALU_DW01_ash_0__n146) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U192 ( .A(ALU_DW01_ash_0__n647), .Y(ALU_DW01_ash_0__n147) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U193 ( .A(ALU_DW01_ash_0__n648), .Y(ALU_DW01_ash_0__n148) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U194 ( .A(ALU_DW01_ash_0__n150), .Y(ALU_DW01_ash_0__n149) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U195 ( .A(ALU_DW01_ash_0__n649), .Y(ALU_DW01_ash_0__n150) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U196 ( .A(ALU_DW01_ash_0__n152), .Y(ALU_DW01_ash_0__n151) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U197 ( .A(ALU_DW01_ash_0__n10), .Y(ALU_DW01_ash_0__n152) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U198 ( .A(ALU_DW01_ash_0__n151), .Y(ALU_DW01_ash_0__n397) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U199 ( .A(ALU_DW01_ash_0__n397), .Y(ALU_DW01_ash_0__n153) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U200 ( .A(ALU_DW01_ash_0__n836), .Y(ALU_DW01_ash_0__n398) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U201 ( .A(ALU_DW01_ash_0__n398), .Y(ALU_DW01_ash_0__n154) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U202 ( .A(ALU_DW01_ash_0__n653), .Y(ALU_DW01_ash_0__n155) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U203 ( .A(ALU_DW01_ash_0__n396), .B(ALU_DW01_ash_0__n650), .Y(ALU_DW01_ash_0__n393) );
  BUFx10_ASAP7_75t_R ALU___ALU_DW01_ash_0___U204 ( .A(ALU_DW01_ash_0__n748), .Y(ALU_DW01_ash_0__n181) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U205 ( .A(ALU_DW01_ash_0__n157), .Y(ALU_DW01_ash_0__n156) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U206 ( .A(ALU_DW01_ash_0__n753), .Y(ALU_DW01_ash_0__n157) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U207 ( .A(ALU_DW01_ash_0__n156), .Y(ALU_DW01_ash_0__n558) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U208 ( .A(ALU_DW01_ash_0__n794), .Y(ALU_DW01_ash_0__n158) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U209 ( .A(ALU_DW01_ash_0__n417), .Y(ALU_DW01_ash_0__n416) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U210 ( .A(ALU_DW01_ash_0__n136), .Y(ALU_DW01_ash_0__n417) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U211 ( .A(ALU_DW01_ash_0__n160), .Y(ALU_DW01_ash_0__n159) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U212 ( .A(ALU_DW01_ash_0__n782), .Y(ALU_DW01_ash_0__n160) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U213 ( .A(ALU_DW01_ash_0__n179), .Y(ALU_DW01_ash_0__n161) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U214 ( .A1(ALU_DW01_ash_0__n663), .A2(ALU_DW01_ash_0__n535), .B1(ALU_DW01_ash_0__n682), .B2(n1068), .C(
        n492), .Y(ALU_DW01_ash_0__n782) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U215 ( .A(ALU_DW01_ash_0__n163), .Y(ALU_DW01_ash_0__n162) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U216 ( .A(ALU_DW01_ash_0__n847), .Y(ALU_DW01_ash_0__n163) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U217 ( .A(ALU_DW01_ash_0__n165), .Y(ALU_DW01_ash_0__n164) );
  AO22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U218 ( .A1(n1064), .A2(ALU_DW01_ash_0__n716), .B1(ALU_DW01_ash_0__n487), .B2(ALU_DW01_ash_0__n702), .Y(
        n793) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U219 ( .A(ALU_DW01_ash_0__n164), .Y(ALU_DW01_ash_0__n506) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U220 ( .A(ALU_DW01_ash_0__n82), .Y(ALU_DW01_ash_0__n167) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U221 ( .A(ALU_DW01_ash_0__n868), .Y(ALU_DW01_ash_0__n168) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U222 ( .A(ALU_DW01_ash_0__n170), .Y(ALU_DW01_ash_0__n169) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U223 ( .A(ALU_DW01_ash_0__n775), .Y(ALU_DW01_ash_0__n170) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U224 ( .A(ALU_DW01_ash_0__n369), .Y(ALU_DW01_ash_0__n664) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U225 ( .A(ALU_DW01_ash_0__n169), .Y(ALU_DW01_ash_0__n594) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U226 ( .A(ALU_DW01_ash_0__n184), .Y(ALU_DW01_ash_0__n171) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U227 ( .A(ALU_DW01_ash_0__n174), .Y(ALU_DW01_ash_0__n172) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U228 ( .A(ALU_DW01_ash_0__n175), .Y(ALU_DW01_ash_0__n173) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U229 ( .A(ALU_DW01_ash_0__n305), .Y(ALU_DW01_ash_0__n174) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U230 ( .A(ALU_DW01_ash_0__n305), .Y(ALU_DW01_ash_0__n175) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U231 ( .A(ALU_DW01_ash_0__n194), .Y(ALU_DW01_ash_0__n176) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U232 ( .A(ALU_DW01_ash_0__n195), .Y(ALU_DW01_ash_0__n194) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U233 ( .A(ALU_DW01_ash_0__n178), .Y(ALU_DW01_ash_0__n177) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U234 ( .A(ALU_DW01_ash_0__n765), .Y(ALU_DW01_ash_0__n178) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U235 ( .A1(ALU_DW01_ash_0__n662), .A2(ALU_DW01_ash_0__n191), .B1(ALU_DW01_ash_0__n681), .B2(n1024), .C(
        n521), .Y(ALU_DW01_ash_0__n765) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U236 ( .A(ALU_DW01_ash_0__n180), .Y(ALU_DW01_ash_0__n179) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U237 ( .A(ALU_DW01_ash_0__n159), .Y(ALU_DW01_ash_0__n180) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U238 ( .A(ALU_DW01_ash_0__n161), .Y(ALU_DW01_ash_0__n491) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U239 ( .A(ALU_DW01_ash_0__n853), .Y(ALU_DW01_ash_0__n598) );
  INVx5_ASAP7_75t_R ALU___ALU_DW01_ash_0___U240 ( .A(ALU_DW01_ash_0__n672), .Y(ALU_DW01_ash_0__n660) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U241 ( .A(ALU_DW01_ash_0__n183), .Y(ALU_DW01_ash_0__n182) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U242 ( .A(ALU_DW01_ash_0__n798), .Y(ALU_DW01_ash_0__n183) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U243 ( .A(ALU_DW01_ash_0__n430), .Y(ALU_DW01_ash_0__n184) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U244 ( .A(ALU_DW01_ash_0__n459), .Y(ALU_DW01_ash_0__n185) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U245 ( .A(ALU_DW01_ash_0__n172), .Y(ALU_DW01_ash_0__n552) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U246 ( .A(ALU_DW01_ash_0__n207), .Y(ALU_DW01_ash_0__n710) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U247 ( .A(ALU_DW01_ash_0__n187), .Y(ALU_DW01_ash_0__n186) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U248 ( .A(ALU_DW01_ash_0__n757), .Y(ALU_DW01_ash_0__n187) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U249 ( .A(ALU_DW01_ash_0__n186), .Y(ALU_DW01_ash_0__n677) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U250 ( .A(ALU_DW01_ash_0__n27), .Y(ALU_DW01_ash_0__n663) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U251 ( .A(ALU_DW01_ash_0__n763), .Y(ALU_DW01_ash_0__n188) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U252 ( .A(ALU_DW01_ash_0__n692), .Y(ALU_DW01_ash_0__n684) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U253 ( .A(ALU_DW01_ash_0__n531), .Y(ALU_DW01_ash_0__n692) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U254 ( .A(ALU_DW01_ash_0__n39), .Y(ALU_DW01_ash_0__n683) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U255 ( .A(n1225), .Y(ALU_DW01_ash_0__n189) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U256 ( .A(n1225), .Y(ALU_DW01_ash_0__n190) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U257 ( .A(n1225), .Y(ALU_DW01_ash_0__n191) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U258 ( .A(n1225), .Y(ALU_DW01_ash_0__n192) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U259 ( .A(ALU_DW01_ash_0__n463), .Y(ALU_DW01_ash_0__n193) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U260 ( .A(ALU_DW01_ash_0__n792), .Y(ALU_DW01_ash_0__n195) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U261 ( .A(ALU_DW01_ash_0__n624), .Y(ALU_DW01_ash_0__n196) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U262 ( .A(ALU_DW01_ash_0__n624), .Y(ALU_DW01_ash_0__n197) );
  CKINVDCx9p33_ASAP7_75t_R ALU___ALU_DW01_ash_0___U263 ( .A(ALU_DW01_ash_0__n176), .Y(ALU_DW01_ash_0__n624) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U264 ( .A(ALU_DW01_ash_0__n199), .Y(ALU_DW01_ash_0__n198) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U265 ( .A(ALU_DW01_ash_0__n828), .Y(ALU_DW01_ash_0__n199) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U266 ( .A(ALU_DW01_ash_0__n607), .B(ALU_DW01_ash_0__n431), .Y(ALU_DW01_ash_0__n828) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U267 ( .A(ALU_DW01_ash_0__n363), .Y(ALU__N267) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U268 ( .A(ALU_DW01_ash_0__n374), .Y(ALU_DW01_ash_0__n201) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U269 ( .A(ALU_DW01_ash_0__n375), .Y(ALU_DW01_ash_0__n202) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U270 ( .A(ALU_DW01_ash_0__n373), .Y(ALU_DW01_ash_0__n203) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U271 ( .A(ALU_DW01_ash_0__n282), .Y(ALU_DW01_ash_0__n204) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U272 ( .A(ALU_DW01_ash_0__n206), .Y(ALU_DW01_ash_0__n205) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U273 ( .A(ALU_DW01_ash_0__n741), .Y(ALU_DW01_ash_0__n206) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U274 ( .A(ALU_DW01_ash_0__n46), .Y(ALU_DW01_ash_0__n207) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U275 ( .A(ALU_DW01_ash_0__n46), .Y(ALU_DW01_ash_0__n208) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U276 ( .A(ALU_DW01_ash_0__n712), .Y(ALU_DW01_ash_0__n209) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U277 ( .A(ALU_DW01_ash_0__n334), .Y(ALU_DW01_ash_0__n712) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U278 ( .A(ALU_DW01_ash_0__n211), .Y(ALU_DW01_ash_0__n210) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U279 ( .A(ALU_DW01_ash_0__n188), .Y(ALU_DW01_ash_0__n211) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U280 ( .A(ALU_DW01_ash_0__n276), .Y(ALU_DW01_ash_0__n584) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U281 ( .A(ALU_DW01_ash_0__n821), .Y(ALU_DW01_ash_0__n212) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U282 ( .A(ALU_DW01_ash_0__n428), .Y(ALU__N266) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U283 ( .A(ALU_DW01_ash_0__n215), .Y(ALU_DW01_ash_0__n214) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U284 ( .A(ALU_DW01_ash_0__n790), .Y(ALU_DW01_ash_0__n215) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U285 ( .A(ALU_DW01_ash_0__n236), .Y(ALU_DW01_ash_0__n216) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U286 ( .A(ALU_DW01_ash_0__n236), .Y(ALU_DW01_ash_0__n217) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U287 ( .A(ALU_DW01_ash_0__n219), .Y(ALU_DW01_ash_0__n218) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U288 ( .A(ALU_DW01_ash_0__n882), .Y(ALU_DW01_ash_0__n219) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U289 ( .A(ALU_DW01_ash_0__n221), .Y(ALU_DW01_ash_0__n220) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U290 ( .A(ALU_DW01_ash_0__n67), .Y(ALU_DW01_ash_0__n221) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U291 ( .A1(n1160), .A2(ALU_DW01_ash_0__n670), .B1(n920), .B2(ALU_DW01_ash_0__n688), .C(
        n455), .Y(ALU_DW01_ash_0__n778) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U292 ( .A(ALU_DW01_ash_0__n223), .Y(ALU_DW01_ash_0__n222) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U293 ( .A(ALU_DW01_ash_0__n127), .Y(ALU_DW01_ash_0__n223) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U294 ( .A(ALU_DW01_ash_0__n308), .Y(ALU_DW01_ash_0__n596) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U295 ( .A(ALU_DW01_ash_0__n225), .Y(ALU_DW01_ash_0__n224) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U296 ( .A(ALU_DW01_ash_0__n761), .Y(ALU_DW01_ash_0__n225) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U297 ( .A1(n1215), .A2(ALU_DW01_ash_0__n666), .B1(ALU_DW01_ash_0__n454), .B2(ALU_DW01_ash_0__n685), .C(
        n384), .Y(ALU_DW01_ash_0__n761) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U298 ( .A(ALU_DW01_ash_0__n227), .Y(ALU_DW01_ash_0__n226) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U299 ( .A(ALU_DW01_ash_0__n806), .Y(ALU_DW01_ash_0__n227) );
  CKINVDCx5p33_ASAP7_75t_R ALU___ALU_DW01_ash_0___U300 ( .A(ALU_DW01_ash_0__n429), .Y(ALU_DW01_ash_0__n571) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U301 ( .A(ALU_DW01_ash_0__n229), .Y(ALU_DW01_ash_0__n228) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U302 ( .A(ALU_DW01_ash_0__n814), .Y(ALU_DW01_ash_0__n229) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U303 ( .A(ALU_DW01_ash_0__n527), .Y(ALU_DW01_ash_0__n665) );
  CKINVDCx5p33_ASAP7_75t_R ALU___ALU_DW01_ash_0___U304 ( .A(ALU_DW01_ash_0__n228), .Y(ALU_DW01_ash_0__n603) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U305 ( .A(ALU_DW01_ash_0__n787), .Y(ALU_DW01_ash_0__n230) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U306 ( .A(ALU_DW01_ash_0__n232), .Y(ALU_DW01_ash_0__n231) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U307 ( .A(ALU_DW01_ash_0__n193), .Y(ALU_DW01_ash_0__n232) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U308 ( .A(ALU_DW01_ash_0__n464), .Y(ALU_DW01_ash_0__n463) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U309 ( .A(ALU_DW01_ash_0__n409), .Y(ALU_DW01_ash_0__n233) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U310 ( .A(ALU_DW01_ash_0__n884), .Y(ALU_DW01_ash_0__n234) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U311 ( .A(ALU_DW01_ash_0__n872), .Y(ALU_DW01_ash_0__n630) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U312 ( .A(ALU_DW01_ash_0__n630), .Y(ALU_DW01_ash_0__n235) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U313 ( .A(ALU_DW01_ash_0__n540), .Y(ALU_DW01_ash_0__n236) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U314 ( .A(ALU_DW01_ash_0__n216), .Y(ALU_DW01_ash_0__n237) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U315 ( .A(ALU_DW01_ash_0__n791), .Y(ALU_DW01_ash_0__n238) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U316 ( .A(ALU_DW01_ash_0__n621), .B(ALU_DW01_ash_0__n185), .Y(ALU_DW01_ash_0__n791) );
  INVx13_ASAP7_75t_R ALU___ALU_DW01_ash_0___U317 ( .A(ALU_DW01_ash_0__n732), .Y(ALU_DW01_ash_0__n621) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U318 ( .A(ALU_DW01_ash_0__n240), .Y(ALU_DW01_ash_0__n239) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U319 ( .A(ALU_DW01_ash_0__n177), .Y(ALU_DW01_ash_0__n240) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U320 ( .A(ALU_DW01_ash_0__n92), .Y(ALU_DW01_ash_0__n520) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U321 ( .A(ALU_DW01_ash_0__n242), .Y(ALU_DW01_ash_0__n241) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U322 ( .A(ALU_DW01_ash_0__n789), .Y(ALU_DW01_ash_0__n242) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U323 ( .A(ALU_DW01_ash_0__n244), .Y(ALU_DW01_ash_0__n243) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U324 ( .A(ALU_DW01_ash_0__n799), .Y(ALU_DW01_ash_0__n244) );
  AO22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U325 ( .A1(ALU_DW01_ash_0__n427), .A2(ALU_DW01_ash_0__n723), .B1(n1060), .B2(ALU_DW01_ash_0__n702), .Y(
        n838) );
  CKINVDCx5p33_ASAP7_75t_R ALU___ALU_DW01_ash_0___U326 ( .A(ALU_DW01_ash_0__n243), .Y(ALU_DW01_ash_0__n580) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U327 ( .A1(ALU_DW01_ash_0__n301), .A2(ALU_DW01_ash_0__n571), .B1(ALU_DW01_ash_0__n413), .B2(ALU_DW01_ash_0__n491), .C(
        n246), .Y(ALU_DW01_ash_0__n864) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U328 ( .A(ALU_DW01_ash_0__n97), .Y(ALU__N279) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U329 ( .A(ALU_DW01_ash_0__n247), .Y(ALU_DW01_ash_0__n246) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U330 ( .A(ALU_DW01_ash_0__n590), .Y(ALU_DW01_ash_0__n247) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U331 ( .A(ALU_DW01_ash_0__n422), .Y(ALU_DW01_ash_0__n731) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U332 ( .A(ALU__n572), .Y(ALU_DW01_ash_0__n248) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U333 ( .A(ALU__n572), .Y(ALU_DW01_ash_0__n249) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U334 ( .A(ALU_DW01_ash_0__n560), .Y(ALU__N265) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U335 ( .A(ALU_DW01_ash_0__n253), .Y(ALU_DW01_ash_0__n251) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U336 ( .A(ALU_DW01_ash_0__n254), .Y(ALU_DW01_ash_0__n252) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U337 ( .A(ALU_DW01_ash_0__n306), .Y(ALU_DW01_ash_0__n253) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U338 ( .A(ALU_DW01_ash_0__n306), .Y(ALU_DW01_ash_0__n254) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U339 ( .A(ALU_DW01_ash_0__n256), .Y(ALU_DW01_ash_0__n255) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U340 ( .A(ALU_DW01_ash_0__n880), .Y(ALU_DW01_ash_0__n256) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U341 ( .A(ALU_DW01_ash_0__n258), .Y(ALU_DW01_ash_0__n257) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U342 ( .A(ALU_DW01_ash_0__n883), .Y(ALU_DW01_ash_0__n258) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U343 ( .A(n1233), .Y(ALU_DW01_ash_0__n259) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U344 ( .A(ALU_DW01_ash_0__n261), .Y(ALU_DW01_ash_0__n260) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U345 ( .A(ALU_DW01_ash_0__n110), .Y(ALU_DW01_ash_0__n261) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U346 ( .A(ALU_DW01_ash_0__n68), .Y(ALU_DW01_ash_0__n477) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U347 ( .A(ALU_DW01_ash_0__n263), .Y(ALU_DW01_ash_0__n262) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U348 ( .A(ALU_DW01_ash_0__n770), .Y(ALU_DW01_ash_0__n263) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U349 ( .A1(n920), .A2(ALU_DW01_ash_0__n670), .B1(n1215), .B2(ALU_DW01_ash_0__n688), .C(
        n586), .Y(ALU_DW01_ash_0__n770) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U350 ( .A(ALU_DW01_ash_0__n265), .Y(ALU_DW01_ash_0__n264) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U351 ( .A(ALU_DW01_ash_0__n766), .Y(ALU_DW01_ash_0__n265) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U352 ( .A(ALU_DW01_ash_0__n264), .Y(ALU_DW01_ash_0__n567) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U353 ( .A(ALU_DW01_ash_0__n803), .Y(ALU_DW01_ash_0__n266) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U354 ( .A1(ALU_DW01_ash_0__n426), .A2(ALU_DW01_ash_0__n446), .B1(ALU_DW01_ash_0__n481), .B2(ALU_DW01_ash_0__n231), .C(
        n268), .Y(ALU_DW01_ash_0__n859) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U355 ( .A(ALU_DW01_ash_0__n61), .Y(ALU__N284) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U356 ( .A(ALU_DW01_ash_0__n269), .Y(ALU_DW01_ash_0__n268) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U357 ( .A(ALU_DW01_ash_0__n797), .Y(ALU_DW01_ash_0__n269) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U358 ( .A(ALU_DW01_ash_0__n320), .Y(ALU__N264) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U359 ( .A(ALU_DW01_ash_0__n780), .Y(ALU_DW01_ash_0__n271) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U360 ( .A(ALU_DW01_ash_0__n767), .Y(ALU_DW01_ash_0__n272) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U361 ( .A1(ALU_DW01_ash_0__n661), .A2(ALU_DW01_ash_0__n487), .B1(ALU_DW01_ash_0__n678), .B2(n1100), .C(
        n474), .Y(ALU_DW01_ash_0__n767) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U362 ( .A(ALU_DW01_ash_0__n348), .Y(ALU_DW01_ash_0__n347) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U363 ( .A(ALU_DW01_ash_0__n103), .Y(ALU_DW01_ash_0__n348) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U364 ( .A(ALU_DW01_ash_0__n772), .Y(ALU_DW01_ash_0__n273) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U365 ( .A(ALU_DW01_ash_0__n275), .Y(ALU_DW01_ash_0__n274) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U366 ( .A(ALU_DW01_ash_0__n783), .Y(ALU_DW01_ash_0__n275) );
  AO221x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U367 ( .A1(ALU_DW01_ash_0__n662), .A2(ALU_DW01_ash_0__n502), .B1(ALU_DW01_ash_0__n679), .B2(n1064), .C(
        n445), .Y(ALU_DW01_ash_0__n783) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U368 ( .A(ALU_DW01_ash_0__n277), .Y(ALU_DW01_ash_0__n276) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U369 ( .A(ALU_DW01_ash_0__n813), .Y(ALU_DW01_ash_0__n277) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U370 ( .A1(ALU_DW01_ash_0__n477), .A2(ALU_DW01_ash_0__n446), .B1(ALU_DW01_ash_0__n599), .B2(ALU_DW01_ash_0__n231), .C(
        n279), .Y(ALU_DW01_ash_0__n861) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U371 ( .A(ALU_DW01_ash_0__n57), .Y(ALU__N282) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U372 ( .A(ALU_DW01_ash_0__n280), .Y(ALU_DW01_ash_0__n279) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U373 ( .A(ALU_DW01_ash_0__n808), .Y(ALU_DW01_ash_0__n280) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U374 ( .A(ALU_DW01_ash_0__n577), .Y(ALU_DW01_ash_0__n281) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U375 ( .A(ALU_DW01_ash_0__n675), .Y(ALU_DW01_ash_0__n662) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U376 ( .A(ALU_DW01_ash_0__n283), .Y(ALU_DW01_ash_0__n730) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U377 ( .A(ALU_DW01_ash_0__n730), .Y(ALU_DW01_ash_0__n282) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U378 ( .A(ALU_DW01_ash_0__n284), .Y(ALU_DW01_ash_0__n283) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U379 ( .A(ALU_DW01_ash_0__n760), .Y(ALU_DW01_ash_0__n284) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U380 ( .A(ALU_DW01_ash_0__n759), .Y(ALU_DW01_ash_0__n285) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U381 ( .A(ALU_DW01_ash_0__n285), .Y(ALU_DW01_ash_0__n333) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U382 ( .A(ALU_DW01_ash_0__n288), .Y(ALU_DW01_ash_0__n286) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U383 ( .A(ALU_DW01_ash_0__n289), .Y(ALU_DW01_ash_0__n287) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U384 ( .A(ALU_DW01_ash_0__n694), .Y(ALU_DW01_ash_0__n288) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U385 ( .A(ALU_DW01_ash_0__n694), .Y(ALU_DW01_ash_0__n289) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U386 ( .A(ALU_DW01_ash_0__n695), .Y(ALU_DW01_ash_0__n694) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U387 ( .A(ALU_DW01_ash_0__n291), .Y(ALU_DW01_ash_0__n290) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U388 ( .A(ALU_DW01_ash_0__n273), .Y(ALU_DW01_ash_0__n291) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U389 ( .A(ALU_DW01_ash_0__n293), .Y(ALU_DW01_ash_0__n292) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U390 ( .A(ALU_DW01_ash_0__n846), .Y(ALU_DW01_ash_0__n293) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U391 ( .A(ALU_DW01_ash_0__n548), .Y(ALU_DW01_ash_0__n294) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U392 ( .A(ALU_DW01_ash_0__n296), .Y(ALU_DW01_ash_0__n295) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U393 ( .A(ALU_DW01_ash_0__n848), .Y(ALU_DW01_ash_0__n296) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U394 ( .A(ALU_DW01_ash_0__n298), .Y(ALU_DW01_ash_0__n297) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U395 ( .A(ALU_DW01_ash_0__n849), .Y(ALU_DW01_ash_0__n298) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U396 ( .A(ALU_DW01_ash_0__n292), .Y(ALU_DW01_ash_0__n548) );
  OR4x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U397 ( .A(ALU_DW01_ash_0__n598), .B(n1164), .C(n352), .D(ALU_DW01_ash_0__n30), .Y(ALU_DW01_ash_0__n846)
         );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U398 ( .A(ALU_DW01_ash_0__n295), .Y(ALU_DW01_ash_0__n549) );
  OR5x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U399 ( .A(ALU_DW01_ash_0__n79), .B(n1123), .C(n1033), .D(ALU_DW01_ash_0__n102), .E(
        n978), .Y(ALU_DW01_ash_0__n848) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U400 ( .A(ALU_DW01_ash_0__n297), .Y(ALU_DW01_ash_0__n550) );
  OR5x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U401 ( .A(ALU_DW01_ash_0__n126), .B(n1208), .C(n619), .D(ALU_DW01_ash_0__n76), .E(ALU_DW01_ash_0__n25), 
        .Y(ALU_DW01_ash_0__n849) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U402 ( .A(ALU_DW01_ash_0__n214), .Y(ALU_DW01_ash_0__n300) );
  CKINVDCx14_ASAP7_75t_R ALU___ALU_DW01_ash_0___U403 ( .A(ALU_DW01_ash_0__n12), .Y(ALU_DW01_ash_0__n619) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U404 ( .A(ALU_DW01_ash_0__n875), .Y(ALU_DW01_ash_0__n588) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U405 ( .A(ALU_DW01_ash_0__n588), .Y(ALU__N268) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U406 ( .A(ALU_DW01_ash_0__n881), .Y(ALU_DW01_ash_0__n501) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U407 ( .A(ALU_DW01_ash_0__n501), .Y(ALU__N262) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U408 ( .A(ALU_DW01_ash_0__n252), .Y(ALU_DW01_ash_0__n304) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U409 ( .A(ALU_DW01_ash_0__n251), .Y(ALU_DW01_ash_0__n305) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U410 ( .A(ALU_DW01_ash_0__n629), .Y(ALU_DW01_ash_0__n306) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U411 ( .A(ALU_DW01_ash_0__n784), .Y(ALU_DW01_ash_0__n307) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U412 ( .A(ALU_DW01_ash_0__n307), .Y(ALU_DW01_ash_0__n629) );
  BUFx10_ASAP7_75t_R ALU___ALU_DW01_ash_0___U413 ( .A(ALU_DW01_ash_0__n810), .Y(ALU_DW01_ash_0__n356) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U414 ( .A(ALU_DW01_ash_0__n309), .Y(ALU_DW01_ash_0__n308) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U415 ( .A(ALU_DW01_ash_0__n809), .Y(ALU_DW01_ash_0__n309) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U416 ( .A(ALU_DW01_ash_0__n262), .Y(ALU_DW01_ash_0__n310) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U417 ( .A(ALU_DW01_ash_0__n855), .Y(ALU__N288) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U418 ( .A1(ALU_DW01_ash_0__n520), .A2(ALU_DW01_ash_0__n611), .B1(ALU_DW01_ash_0__n567), .B2(ALU_DW01_ash_0__n618), .C1(
        n473), .C2(ALU_DW01_ash_0__n461), .Y(ALU_DW01_ash_0__n764) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U419 ( .A(ALU_DW01_ash_0__n137), .Y(ALU_DW01_ash_0__n312) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U420 ( .A1(ALU_DW01_ash_0__n411), .A2(ALU_DW01_ash_0__n591), .B1(ALU_DW01_ash_0__n312), .B2(ALU_DW01_ash_0__n626), .Y(
        n762) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U421 ( .A(ALU_DW01_ash_0__n138), .Y(ALU_DW01_ash_0__n313) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U422 ( .A(ALU_DW01_ash_0__n347), .Y(ALU_DW01_ash_0__n473) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U423 ( .A1(ALU_DW01_ash_0__n580), .A2(ALU_DW01_ash_0__n619), .B1(ALU_DW01_ash_0__n594), .B2(ALU_DW01_ash_0__n331), .C(
        n315), .Y(ALU_DW01_ash_0__n867) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U424 ( .A(ALU_DW01_ash_0__n98), .Y(ALU__N276) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U425 ( .A(ALU_DW01_ash_0__n316), .Y(ALU_DW01_ash_0__n315) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U426 ( .A(ALU_DW01_ash_0__n825), .Y(ALU_DW01_ash_0__n316) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U427 ( .A(ALU_DW01_ash_0__n675), .Y(ALU_DW01_ash_0__n317) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U428 ( .A(ALU_DW01_ash_0__n29), .Y(ALU_DW01_ash_0__n318) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U429 ( .A(n858), .Y(ALU_DW01_ash_0__n319) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U430 ( .A(ALU_DW01_ash_0__n879), .Y(ALU_DW01_ash_0__n608) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U431 ( .A(ALU_DW01_ash_0__n608), .Y(ALU_DW01_ash_0__n320) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U432 ( .A(ALU_DW01_ash_0__n727), .Y(ALU_DW01_ash_0__n321) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U433 ( .A(ALU_DW01_ash_0__n727), .Y(ALU_DW01_ash_0__n322) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U434 ( .A(ALU_DW01_ash_0__n727), .Y(ALU_DW01_ash_0__n323) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U435 ( .A(ALU_DW01_ash_0__n727), .Y(ALU_DW01_ash_0__n324) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U436 ( .A(ALU_DW01_ash_0__n323), .Y(ALU_DW01_ash_0__n726) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U437 ( .A(ALU_DW01_ash_0__n372), .Y(ALU_DW01_ash_0__n727) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U438 ( .A(ALU_DW01_ash_0__n750), .Y(ALU_DW01_ash_0__n325) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U439 ( .A(ALU_DW01_ash_0__n327), .Y(ALU_DW01_ash_0__n326) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U440 ( .A(ALU_DW01_ash_0__n747), .Y(ALU_DW01_ash_0__n327) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U441 ( .A(ALU_DW01_ash_0__n329), .Y(ALU_DW01_ash_0__n328) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U442 ( .A(ALU_DW01_ash_0__n786), .Y(ALU_DW01_ash_0__n329) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U443 ( .A(ALU_DW01_ash_0__n546), .Y(ALU_DW01_ash_0__n330) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U444 ( .A(ALU_DW01_ash_0__n546), .Y(ALU_DW01_ash_0__n331) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U445 ( .A(ALU_DW01_ash_0__n546), .Y(ALU_DW01_ash_0__n332) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U446 ( .A(ALU_DW01_ash_0__n286), .Y(ALU_DW01_ash_0__n689) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U447 ( .A(ALU_DW01_ash_0__n287), .Y(ALU_DW01_ash_0__n532) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U448 ( .A(ALU_DW01_ash_0__n340), .B(ALU_DW01_ash_0__n631), .Y(ALU_DW01_ash_0__n759) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U449 ( .A(ALU_DW01_ash_0__n713), .Y(ALU_DW01_ash_0__n334) );
  INVx5_ASAP7_75t_R ALU___ALU_DW01_ash_0___U450 ( .A(ALU_DW01_ash_0__n333), .Y(ALU_DW01_ash_0__n713) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U451 ( .A(ALU_DW01_ash_0__n336), .Y(ALU_DW01_ash_0__n335) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U452 ( .A(ALU_DW01_ash_0__n271), .Y(ALU_DW01_ash_0__n336) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U453 ( .A1(ALU_DW01_ash_0__n473), .A2(ALU_DW01_ash_0__n446), .B1(ALU_DW01_ash_0__n416), .B2(ALU_DW01_ash_0__n231), .C(
        n338), .Y(ALU_DW01_ash_0__n858) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U454 ( .A(ALU_DW01_ash_0__n48), .Y(ALU__N285) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U455 ( .A(ALU_DW01_ash_0__n339), .Y(ALU_DW01_ash_0__n338) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U456 ( .A(ALU_DW01_ash_0__n795), .Y(ALU_DW01_ash_0__n339) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U457 ( .A(ALU_DW01_ash_0__n494), .Y(ALU_DW01_ash_0__n341) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U458 ( .A(ALU_DW01_ash_0__n494), .Y(ALU_DW01_ash_0__n342) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U459 ( .A(ALU_DW01_ash_0__n494), .Y(ALU_DW01_ash_0__n343) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U460 ( .A(ALU_DW01_ash_0__n458), .Y(ALU_DW01_ash_0__n344) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U461 ( .A(ALU_DW01_ash_0__n459), .Y(ALU_DW01_ash_0__n458) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U462 ( .A(ALU_DW01_ash_0__n386), .Y(ALU_DW01_ash_0__n345) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U463 ( .A(ALU_DW01_ash_0__n386), .Y(ALU_DW01_ash_0__n346) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U464 ( .A(ALU_DW01_ash_0__n528), .Y(ALU_DW01_ash_0__n661) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U465 ( .A(ALU_DW01_ash_0__n350), .Y(ALU_DW01_ash_0__n349) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U466 ( .A(ALU_DW01_ash_0__n88), .Y(ALU_DW01_ash_0__n350) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U467 ( .A(ALU_DW01_ash_0__n526), .Y(ALU_DW01_ash_0__n667) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U468 ( .A(ALU_DW01_ash_0__n51), .Y(ALU_DW01_ash_0__n509) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U469 ( .A(ALU_DW01_ash_0__n829), .Y(ALU_DW01_ash_0__n351) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U470 ( .A(ALU_DW01_ash_0__n635), .B(ALU_DW01_ash_0__n636), .Y(ALU_DW01_ash_0__n352) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U471 ( .A(ALU_DW01_ash_0__n660), .B(n925), .Y(ALU_DW01_ash_0__n633) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U472 ( .A(ALU_DW01_ash_0__n132), .Y(ALU_DW01_ash_0__n353) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U473 ( .A(ALU_DW01_ash_0__n683), .B(n1073), .Y(ALU_DW01_ash_0__n634) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U474 ( .A(ALU_DW01_ash_0__n133), .Y(ALU_DW01_ash_0__n354) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U475 ( .A(ALU_DW01_ash_0__n353), .B(ALU_DW01_ash_0__n354), .Y(ALU_DW01_ash_0__n637) );
  OR3x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U476 ( .A(ALU_DW01_ash_0__n621), .B(ALU_DW01_ash_0__n472), .C(ALU_DW01_ash_0__n601), .Y(ALU_DW01_ash_0__n880) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U477 ( .A(ALU_DW01_ash_0__n255), .Y(ALU__N263) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U478 ( .A1(ALU_DW01_ash_0__n520), .A2(ALU_DW01_ash_0__n414), .B1(ALU_DW01_ash_0__n388), .B2(ALU_DW01_ash_0__n193), .C(
        n359), .Y(ALU_DW01_ash_0__n862) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U479 ( .A(ALU_DW01_ash_0__n63), .Y(ALU__N281) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U480 ( .A(ALU_DW01_ash_0__n360), .Y(ALU_DW01_ash_0__n359) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U481 ( .A(ALU_DW01_ash_0__n812), .Y(ALU_DW01_ash_0__n360) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U482 ( .A(ALU_DW01_ash_0__n529), .Y(ALU__N274) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U483 ( .A(ALU_DW01_ash_0__n556), .Y(ALU__N272) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U484 ( .A(ALU_DW01_ash_0__n876), .Y(ALU_DW01_ash_0__n614) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U485 ( .A(ALU_DW01_ash_0__n614), .Y(ALU_DW01_ash_0__n363) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U486 ( .A(ALU__n731), .Y(ALU_DW01_ash_0__n364) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U487 ( .A(ALU_DW01_ash_0__n616), .Y(ALU_DW01_ash_0__n679) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U488 ( .A(ALU_DW01_ash_0__n289), .Y(ALU_DW01_ash_0__n616) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U489 ( .A(ALU_DW01_ash_0__n366), .Y(ALU_DW01_ash_0__n365) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U490 ( .A(ALU_DW01_ash_0__n205), .Y(ALU_DW01_ash_0__n366) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U491 ( .A(ALU_DW01_ash_0__n746), .Y(ALU_DW01_ash_0__n367) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U492 ( .A(ALU_DW01_ash_0__n370), .Y(ALU_DW01_ash_0__n368) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U493 ( .A(ALU_DW01_ash_0__n371), .Y(ALU_DW01_ash_0__n369) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U494 ( .A(ALU_DW01_ash_0__n45), .Y(ALU_DW01_ash_0__n370) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U495 ( .A(ALU_DW01_ash_0__n44), .Y(ALU_DW01_ash_0__n371) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U496 ( .A(ALU_DW01_ash_0__n35), .Y(ALU_DW01_ash_0__n672) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U497 ( .A(ALU_DW01_ash_0__n317), .Y(ALU_DW01_ash_0__n674) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U498 ( .A(ALU_DW01_ash_0__n374), .Y(ALU_DW01_ash_0__n372) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U499 ( .A(ALU_DW01_ash_0__n375), .Y(ALU_DW01_ash_0__n373) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U500 ( .A(ALU_DW01_ash_0__n65), .Y(ALU_DW01_ash_0__n374) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U501 ( .A(ALU_DW01_ash_0__n49), .Y(ALU_DW01_ash_0__n375) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U502 ( .A(ALU_DW01_ash_0__n373), .Y(ALU_DW01_ash_0__n728) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U503 ( .A(ALU_DW01_ash_0__n282), .Y(ALU_DW01_ash_0__n729) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U504 ( .A(ALU_DW01_ash_0__n66), .Y(ALU_DW01_ash_0__n376) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U505 ( .A(ALU_DW01_ash_0__n709), .Y(ALU_DW01_ash_0__n377) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U506 ( .A(ALU_DW01_ash_0__n209), .Y(ALU_DW01_ash_0__n706) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U507 ( .A(ALU_DW01_ash_0__n711), .Y(ALU_DW01_ash_0__n709) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U508 ( .A(ALU_DW01_ash_0__n379), .Y(ALU_DW01_ash_0__n378) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U509 ( .A(ALU_DW01_ash_0__n328), .Y(ALU_DW01_ash_0__n379) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U510 ( .A(ALU_DW01_ash_0__n617), .Y(ALU_DW01_ash_0__n380) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U511 ( .A1(ALU_DW01_ash_0__n603), .A2(ALU_DW01_ash_0__n619), .B1(ALU_DW01_ash_0__n567), .B2(ALU_DW01_ash_0__n330), .C(
        n382), .Y(ALU_DW01_ash_0__n866) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U512 ( .A(ALU_DW01_ash_0__n87), .Y(ALU__N277) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U513 ( .A(ALU_DW01_ash_0__n383), .Y(ALU_DW01_ash_0__n382) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U514 ( .A(ALU_DW01_ash_0__n823), .Y(ALU_DW01_ash_0__n383) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U515 ( .A(ALU_DW01_ash_0__n768), .Y(ALU_DW01_ash_0__n384) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U516 ( .A(ALU_DW01_ash_0__n346), .Y(ALU_DW01_ash_0__n385) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U517 ( .A(ALU_DW01_ash_0__n613), .Y(ALU_DW01_ash_0__n386) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U518 ( .A(ALU_DW01_ash_0__n752), .Y(ALU_DW01_ash_0__n387) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U519 ( .A(ALU_DW01_ash_0__n391), .Y(ALU_DW01_ash_0__n390) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U520 ( .A(ALU_DW01_ash_0__n274), .Y(ALU_DW01_ash_0__n391) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U521 ( .A(n1091), .Y(ALU_DW01_ash_0__n392) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U522 ( .A(ALU_DW01_ash_0__n666), .B(n929), .Y(ALU_DW01_ash_0__n647) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U523 ( .A(ALU_DW01_ash_0__n147), .Y(ALU_DW01_ash_0__n394) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U524 ( .A(ALU_DW01_ash_0__n683), .B(n1029), .Y(ALU_DW01_ash_0__n648) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U525 ( .A(ALU_DW01_ash_0__n148), .Y(ALU_DW01_ash_0__n395) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U526 ( .A(ALU_DW01_ash_0__n154), .Y(ALU_DW01_ash_0__n649) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U527 ( .A(ALU_DW01_ash_0__n149), .Y(ALU_DW01_ash_0__n396) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U528 ( .A(ALU_DW01_ash_0__n394), .B(ALU_DW01_ash_0__n395), .Y(ALU_DW01_ash_0__n651) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U529 ( .A(ALU_DW01_ash_0__n400), .B(ALU_DW01_ash_0__n399), .Y(ALU_DW01_ash_0__n836) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U530 ( .A(n973), .B(ALU_DW01_ash_0__n722), .Y(ALU_DW01_ash_0__n653) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U531 ( .A(ALU_DW01_ash_0__n155), .Y(ALU_DW01_ash_0__n399) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U532 ( .A(ALU_DW01_ash_0__n553), .B(ALU_DW01_ash_0__n702), .Y(ALU_DW01_ash_0__n652) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U533 ( .A(ALU_DW01_ash_0__n652), .Y(ALU_DW01_ash_0__n400) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U534 ( .A(ALU_DW01_ash_0__n21), .Y(ALU_DW01_ash_0__n743) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U535 ( .A(ALU_DW01_ash_0__n16), .Y(ALU_DW01_ash_0__n401) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U536 ( .A(ALU_DW01_ash_0__n533), .B(ALU_DW01_ash_0__n669), .Y(ALU_DW01_ash_0__n655) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U537 ( .A(ALU_DW01_ash_0__n655), .Y(ALU_DW01_ash_0__n402) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U538 ( .A(n1060), .B(ALU_DW01_ash_0__n33), .Y(ALU_DW01_ash_0__n656) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U539 ( .A(ALU_DW01_ash_0__n17), .Y(ALU_DW01_ash_0__n403) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U540 ( .A(ALU_DW01_ash_0__n406), .B(ALU_DW01_ash_0__n407), .Y(ALU_DW01_ash_0__n404) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U541 ( .A(ALU_DW01_ash_0__n18), .B(ALU_DW01_ash_0__n22), .Y(ALU_DW01_ash_0__n654) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U542 ( .A(ALU_DW01_ash_0__n402), .B(ALU_DW01_ash_0__n403), .Y(ALU_DW01_ash_0__n657) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U543 ( .A(n964), .B(ALU_DW01_ash_0__n726), .Y(ALU_DW01_ash_0__n658) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U544 ( .A(ALU_DW01_ash_0__n23), .Y(ALU_DW01_ash_0__n406) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U545 ( .A(n1015), .B(ALU_DW01_ash_0__n706), .Y(ALU_DW01_ash_0__n659) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U546 ( .A(ALU_DW01_ash_0__n24), .Y(ALU_DW01_ash_0__n407) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U547 ( .A(ALU__n503), .Y(ALU_DW01_ash_0__n408) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U548 ( .A(ALU__n503), .Y(ALU_DW01_ash_0__n409) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U549 ( .A(ALU__n503), .Y(ALU_DW01_ash_0__n410) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U550 ( .A(ALU__n503), .Y(ALU_DW01_ash_0__n411) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_ash_0___U551 ( .A(ALU_DW01_ash_0__n818), .Y(ALU_DW01_ash_0__n412) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U552 ( .A(ALU_DW01_ash_0__n448), .Y(ALU_DW01_ash_0__n413) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U553 ( .A(ALU_DW01_ash_0__n448), .Y(ALU_DW01_ash_0__n414) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U554 ( .A(ALU__n794), .Y(ALU_DW01_ash_0__n415) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U555 ( .A(ALU_DW01_ash_0__n419), .Y(ALU_DW01_ash_0__n418) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U556 ( .A(ALU_DW01_ash_0__n800), .Y(ALU_DW01_ash_0__n419) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U557 ( .A(ALU_DW01_ash_0__n418), .Y(ALU_DW01_ash_0__n564) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U558 ( .A1(ALU_DW01_ash_0__n477), .A2(ALU_DW01_ash_0__n611), .B1(ALU_DW01_ash_0__n558), .B2(ALU_DW01_ash_0__n618), .C1(
        n506), .C2(ALU_DW01_ash_0__n462), .Y(ALU_DW01_ash_0__n750) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U559 ( .A(ALU_DW01_ash_0__n325), .Y(ALU_DW01_ash_0__n420) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U560 ( .A1(ALU_DW01_ash_0__n410), .A2(ALU_DW01_ash_0__n517), .B1(ALU_DW01_ash_0__n420), .B2(ALU_DW01_ash_0__n626), .Y(
        n747) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U561 ( .A(ALU_DW01_ash_0__n326), .Y(ALU_DW01_ash_0__n421) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_ash_0___U562 ( .A(ALU_DW01_ash_0__n423), .Y(ALU_DW01_ash_0__n422) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_ash_0___U563 ( .A(ALU_DW01_ash_0__n412), .Y(ALU_DW01_ash_0__n423) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U564 ( .A(ALU_DW01_ash_0__n425), .Y(ALU_DW01_ash_0__n424) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U565 ( .A(ALU_DW01_ash_0__n801), .Y(ALU_DW01_ash_0__n425) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U566 ( .A(ALU_DW01_ash_0__n534), .Y(ALU_DW01_ash_0__n427) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U567 ( .A(ALU_DW01_ash_0__n877), .Y(ALU_DW01_ash_0__n620) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U568 ( .A(ALU_DW01_ash_0__n620), .Y(ALU_DW01_ash_0__n428) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U569 ( .A(ALU_DW01_ash_0__n226), .Y(ALU_DW01_ash_0__n429) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U570 ( .A(ALU_DW01_ash_0__n431), .Y(ALU_DW01_ash_0__n430) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U571 ( .A(ALU_DW01_ash_0__n432), .Y(ALU_DW01_ash_0__n431) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U572 ( .A(ALU_DW01_ash_0__n472), .Y(ALU_DW01_ash_0__n432) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U573 ( .A(ALU__n901), .Y(ALU_DW01_ash_0__n472) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U574 ( .A(ALU_DW01_ash_0__n665), .B(ALU_DW01_ash_0__n47), .Y(ALU_DW01_ash_0__n640) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U575 ( .A(ALU_DW01_ash_0__n117), .Y(ALU_DW01_ash_0__n434) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U576 ( .A(ALU_DW01_ash_0__n683), .B(n969), .Y(ALU_DW01_ash_0__n641) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U577 ( .A(ALU_DW01_ash_0__n118), .Y(ALU_DW01_ash_0__n435) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U578 ( .A(ALU_DW01_ash_0__n124), .Y(ALU_DW01_ash_0__n642) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U579 ( .A(ALU_DW01_ash_0__n119), .Y(ALU_DW01_ash_0__n436) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U580 ( .A(ALU_DW01_ash_0__n434), .B(ALU_DW01_ash_0__n435), .Y(ALU_DW01_ash_0__n644) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U581 ( .A(ALU_DW01_ash_0__n439), .B(ALU_DW01_ash_0__n440), .Y(ALU_DW01_ash_0__n834) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U582 ( .A(ALU_DW01_ash_0__n142), .B(ALU_DW01_ash_0__n702), .Y(ALU_DW01_ash_0__n645) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U583 ( .A(ALU_DW01_ash_0__n125), .Y(ALU_DW01_ash_0__n439) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U584 ( .A(ALU_DW01_ash_0__n281), .B(ALU_DW01_ash_0__n722), .Y(ALU_DW01_ash_0__n646) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U585 ( .A(ALU_DW01_ash_0__n646), .Y(ALU_DW01_ash_0__n440) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U586 ( .A(ALU_DW01_ash_0__n42), .Y(ALU_DW01_ash_0__n722) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U587 ( .A1(ALU_DW01_ash_0__n506), .A2(ALU_DW01_ash_0__n547), .B1(ALU_DW01_ash_0__n378), .B2(ALU_DW01_ash_0__n230), .C(
        n442), .Y(ALU_DW01_ash_0__n857) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U588 ( .A(ALU_DW01_ash_0__n41), .Y(ALU__N286) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U589 ( .A(ALU_DW01_ash_0__n443), .Y(ALU_DW01_ash_0__n442) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U590 ( .A(ALU_DW01_ash_0__n788), .Y(ALU_DW01_ash_0__n443) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U591 ( .A(ALU_DW01_ash_0__n390), .Y(ALU_DW01_ash_0__n444) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U592 ( .A(ALU_DW01_ash_0__n807), .Y(ALU_DW01_ash_0__n445) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U593 ( .A(ALU_DW01_ash_0__n414), .Y(ALU_DW01_ash_0__n446) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U594 ( .A(ALU_DW01_ash_0__n413), .Y(ALU_DW01_ash_0__n447) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U595 ( .A(ALU_DW01_ash_0__n547), .Y(ALU_DW01_ash_0__n448) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U596 ( .A(ALU_DW01_ash_0__n744), .Y(ALU_DW01_ash_0__n449) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U597 ( .A(ALU_DW01_ash_0__n451), .Y(ALU_DW01_ash_0__n450) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U598 ( .A(ALU_DW01_ash_0__n198), .Y(ALU_DW01_ash_0__n451) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U599 ( .A(ALU_DW01_ash_0__n453), .Y(ALU_DW01_ash_0__n452) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U600 ( .A(ALU_DW01_ash_0__n769), .Y(ALU_DW01_ash_0__n453) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U601 ( .A(n1010), .Y(ALU_DW01_ash_0__n454) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U602 ( .A(ALU_DW01_ash_0__n785), .Y(ALU_DW01_ash_0__n455) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U603 ( .A(ALU_DW01_ash_0__n220), .Y(ALU_DW01_ash_0__n456) );
  AO22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U604 ( .A1(ALU_DW01_ash_0__n706), .A2(n1100), .B1(ALU_DW01_ash_0__n715), .B2(ALU_DW01_ash_0__n487), .Y(
        n785) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U605 ( .A(n1174), .Y(ALU_DW01_ash_0__n457) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U606 ( .A(ALU_DW01_ash_0__n756), .Y(ALU_DW01_ash_0__n459) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U607 ( .A(ALU_DW01_ash_0__n625), .Y(ALU_DW01_ash_0__n460) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U608 ( .A(ALU_DW01_ash_0__n625), .Y(ALU_DW01_ash_0__n461) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U609 ( .A(ALU_DW01_ash_0__n625), .Y(ALU_DW01_ash_0__n462) );
  CKINVDCx8_ASAP7_75t_R ALU___ALU_DW01_ash_0___U610 ( .A(ALU_DW01_ash_0__n171), .Y(ALU_DW01_ash_0__n735) );
  CKINVDCx14_ASAP7_75t_R ALU___ALU_DW01_ash_0___U611 ( .A(ALU_DW01_ash_0__n344), .Y(ALU_DW01_ash_0__n625) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U612 ( .A(ALU_DW01_ash_0__n230), .Y(ALU_DW01_ash_0__n464) );
  OR2x4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U613 ( .A(ALU_DW01_ash_0__n626), .B(ALU_DW01_ash_0__n551), .Y(ALU_DW01_ash_0__n787) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U614 ( .A(ALU_DW01_ash_0__n466), .Y(ALU_DW01_ash_0__n465) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U615 ( .A(ALU_DW01_ash_0__n874), .Y(ALU_DW01_ash_0__n466) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U616 ( .A1(ALU_DW01_ash_0__n509), .A2(ALU_DW01_ash_0__n611), .B1(ALU_DW01_ash_0__n594), .B2(ALU_DW01_ash_0__n618), .C1(
        n426), .C2(ALU_DW01_ash_0__n462), .Y(ALU_DW01_ash_0__n773) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U617 ( .A(ALU_DW01_ash_0__n107), .Y(ALU_DW01_ash_0__n467) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U618 ( .A1(ALU_DW01_ash_0__n233), .A2(ALU_DW01_ash_0__n543), .B1(ALU_DW01_ash_0__n467), .B2(ALU_DW01_ash_0__n626), .Y(
        n771) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U619 ( .A(ALU_DW01_ash_0__n108), .Y(ALU_DW01_ash_0__n468) );
  O2A1O1Ixp33_ASAP7_75t_R ALU___ALU_DW01_ash_0___U620 ( .A1(ALU_DW01_ash_0__n310), .A2(ALU_DW01_ash_0__n367), .B(ALU_DW01_ash_0__n468), .C(ALU_DW01_ash_0__n551), .Y(
        n855) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U621 ( .A1(ALU_DW01_ash_0__n444), .A2(ALU_DW01_ash_0__n449), .B1(ALU_DW01_ash_0__n575), .B2(ALU_DW01_ash_0__n464), .C(
        n470), .Y(ALU_DW01_ash_0__n860) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U622 ( .A(ALU_DW01_ash_0__n52), .Y(ALU__N283) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U623 ( .A(ALU_DW01_ash_0__n471), .Y(ALU_DW01_ash_0__n470) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U624 ( .A(ALU_DW01_ash_0__n802), .Y(ALU_DW01_ash_0__n471) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U625 ( .A(ALU_DW01_ash_0__n796), .Y(ALU_DW01_ash_0__n474) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U626 ( .A1(ALU_DW01_ash_0__n503), .A2(ALU_DW01_ash_0__n716), .B1(n1064), .B2(ALU_DW01_ash_0__n702), .Y(
        n796) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U627 ( .A(ALU_DW01_ash_0__n476), .Y(ALU_DW01_ash_0__n475) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U628 ( .A(ALU_DW01_ash_0__n811), .Y(ALU_DW01_ash_0__n476) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U629 ( .A(ALU_DW01_ash_0__n869), .Y(ALU_DW01_ash_0__n478) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U630 ( .A(ALU_DW01_ash_0__n480), .Y(ALU_DW01_ash_0__n479) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U631 ( .A(ALU_DW01_ash_0__n873), .Y(ALU_DW01_ash_0__n480) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U632 ( .A(ALU_DW01_ash_0__n690), .Y(ALU_DW01_ash_0__n682) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U633 ( .A(ALU_DW01_ash_0__n531), .Y(ALU_DW01_ash_0__n690) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U634 ( .A(ALU_DW01_ash_0__n622), .B(ALU_DW01_ash_0__n447), .Y(ALU_DW01_ash_0__n882) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U635 ( .A(ALU_DW01_ash_0__n218), .Y(ALU__N261) );
  OR5x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U636 ( .A(ALU_DW01_ash_0__n485), .B(n1162), .C(n1075), .D(n701), .E(
        n415), .Y(ALU_DW01_ash_0__n847) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U637 ( .A(ALU_DW01_ash_0__n162), .Y(ALU_DW01_ash_0__n484) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U638 ( .A(ALU_DW01_ash_0__n852), .Y(ALU_DW01_ash_0__n485) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U639 ( .A(ALU__n936), .Y(ALU_DW01_ash_0__n486) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U640 ( .A(ALU__n936), .Y(ALU_DW01_ash_0__n487) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U641 ( .A1(ALU_DW01_ash_0__n565), .A2(ALU_DW01_ash_0__n619), .B1(ALU_DW01_ash_0__n558), .B2(ALU_DW01_ash_0__n330), .C(
        n489), .Y(ALU_DW01_ash_0__n865) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U642 ( .A(ALU_DW01_ash_0__n77), .Y(ALU__N278) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U643 ( .A(ALU_DW01_ash_0__n490), .Y(ALU_DW01_ash_0__n489) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U644 ( .A(ALU_DW01_ash_0__n820), .Y(ALU_DW01_ash_0__n490) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U645 ( .A(ALU_DW01_ash_0__n432), .B(ALU_DW01_ash_0__n248), .Y(ALU_DW01_ash_0__n784) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U646 ( .A(ALU_DW01_ash_0__n551), .B(ALU_DW01_ash_0__n411), .Y(ALU_DW01_ash_0__n830) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U647 ( .A(ALU_DW01_ash_0__n819), .Y(ALU_DW01_ash_0__n492) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U648 ( .A(ALU_DW01_ash_0__n871), .Y(ALU_DW01_ash_0__n493) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U649 ( .A(n892), .Y(ALU_DW01_ash_0__n494) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U650 ( .A(ALU_DW01_ash_0__n496), .Y(ALU_DW01_ash_0__n495) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U651 ( .A(ALU_DW01_ash_0__n452), .Y(ALU_DW01_ash_0__n496) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U652 ( .A(ALU_DW01_ash_0__n495), .Y(ALU_DW01_ash_0__n622) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U653 ( .A(ALU_DW01_ash_0__n378), .B(ALU_DW01_ash_0__n621), .Y(ALU_DW01_ash_0__n873) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U654 ( .A(ALU_DW01_ash_0__n479), .Y(ALU__N270) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U655 ( .A(ALU_DW01_ash_0__n564), .B(ALU_DW01_ash_0__n447), .Y(ALU_DW01_ash_0__n883) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U656 ( .A(ALU_DW01_ash_0__n257), .Y(ALU__N260) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U657 ( .A(ALU_DW01_ash_0__n758), .Y(ALU_DW01_ash_0__n499) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U658 ( .A(ALU_DW01_ash_0__n105), .Y(ALU_DW01_ash_0__n500) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U659 ( .A(ALU_DW01_ash_0__n401), .B(ALU_DW01_ash_0__n446), .Y(ALU_DW01_ash_0__n881) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U660 ( .A(n1178), .Y(ALU_DW01_ash_0__n502) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U661 ( .A(n1178), .Y(ALU_DW01_ash_0__n503) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U662 ( .A(ALU__n968), .Y(ALU_DW01_ash_0__n504) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U663 ( .A(ALU_DW01_ash_0__n793), .Y(ALU_DW01_ash_0__n505) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U664 ( .A(ALU_DW01_ash_0__n249), .Y(ALU_DW01_ash_0__n507) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U665 ( .A(ALU_DW01_ash_0__n248), .Y(ALU_DW01_ash_0__n508) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U666 ( .A(ALU_DW01_ash_0__n817), .Y(ALU_DW01_ash_0__n510) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U667 ( .A(ALU_DW01_ash_0__n692), .Y(ALU_DW01_ash_0__n615) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U668 ( .A(ALU_DW01_ash_0__n416), .B(ALU_DW01_ash_0__n621), .Y(ALU_DW01_ash_0__n874) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U669 ( .A(ALU_DW01_ash_0__n465), .Y(ALU__N269) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U670 ( .A(ALU_DW01_ash_0__n856), .Y(ALU__N287) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U671 ( .A(ALU_DW01_ash_0__n779), .Y(ALU_DW01_ash_0__n513) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U672 ( .A1(ALU_DW01_ash_0__n509), .A2(ALU_DW01_ash_0__n332), .B1(ALU_DW01_ash_0__n365), .B2(ALU_DW01_ash_0__n232), .C(
        n515), .Y(ALU_DW01_ash_0__n863) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U673 ( .A(ALU_DW01_ash_0__n70), .Y(ALU__N280) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U674 ( .A(ALU_DW01_ash_0__n516), .Y(ALU_DW01_ash_0__n515) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U675 ( .A(ALU_DW01_ash_0__n816), .Y(ALU_DW01_ash_0__n516) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U676 ( .A1(ALU_DW01_ash_0__n380), .A2(ALU_DW01_ash_0__n401), .B1(ALU_DW01_ash_0__n385), .B2(ALU_DW01_ash_0__n565), .C(
        n518), .Y(ALU_DW01_ash_0__n749) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U677 ( .A(ALU_DW01_ash_0__n222), .Y(ALU_DW01_ash_0__n517) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U678 ( .A(ALU_DW01_ash_0__n519), .Y(ALU_DW01_ash_0__n518) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U679 ( .A(ALU_DW01_ash_0__n831), .Y(ALU_DW01_ash_0__n519) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U680 ( .A(ALU_DW01_ash_0__n815), .Y(ALU_DW01_ash_0__n521) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U681 ( .A(ALU_DW01_ash_0__n40), .Y(ALU_DW01_ash_0__n681) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U682 ( .A(ALU_DW01_ash_0__n839), .Y(ALU_DW01_ash_0__n523) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U683 ( .A(ALU_DW01_ash_0__n525), .Y(ALU_DW01_ash_0__n524) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U684 ( .A(ALU_DW01_ash_0__n234), .Y(ALU_DW01_ash_0__n525) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U685 ( .A(ALU_DW01_ash_0__n208), .Y(ALU_DW01_ash_0__n711) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U686 ( .A(ALU_DW01_ash_0__n34), .Y(ALU_DW01_ash_0__n526) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U687 ( .A(ALU_DW01_ash_0__n26), .Y(ALU_DW01_ash_0__n527) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U688 ( .A(ALU_DW01_ash_0__n527), .Y(ALU_DW01_ash_0__n666) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U689 ( .A(ALU_DW01_ash_0__n526), .Y(ALU_DW01_ash_0__n668) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U690 ( .A(ALU_DW01_ash_0__n530), .Y(ALU_DW01_ash_0__n529) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U691 ( .A(ALU_DW01_ash_0__n478), .Y(ALU_DW01_ash_0__n530) );
  CKINVDCx12_ASAP7_75t_R ALU___ALU_DW01_ash_0___U692 ( .A(ALU_DW01_ash_0__n687), .Y(ALU_DW01_ash_0__n531) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U693 ( .A(ALU__n905), .Y(ALU_DW01_ash_0__n533) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U694 ( .A(ALU__n905), .Y(ALU_DW01_ash_0__n534) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U695 ( .A(ALU__n904), .Y(ALU_DW01_ash_0__n535) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U696 ( .A(ALU__n904), .Y(ALU_DW01_ash_0__n536) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U697 ( .A(ALU__n904), .Y(ALU_DW01_ash_0__n537) );
  AO22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U698 ( .A1(ALU_DW01_ash_0__n537), .A2(ALU_DW01_ash_0__n717), .B1(n1068), .B2(ALU_DW01_ash_0__n698), .Y(
        n815) );
  AO22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U699 ( .A1(n1182), .A2(ALU_DW01_ash_0__n718), .B1(ALU_DW01_ash_0__n536), .B2(ALU_DW01_ash_0__n699), .Y(
        n817) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U700 ( .A(n749), .B(ALU_DW01_ash_0__n341), .Y(ALU_DW01_ash_0__n623) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U701 ( .A(ALU_DW01_ash_0__n237), .Y(ALU_DW01_ash_0__n538) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U702 ( .A(ALU_DW01_ash_0__n217), .Y(ALU_DW01_ash_0__n539) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U703 ( .A(ALU_DW01_ash_0__n238), .Y(ALU_DW01_ash_0__n540) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U704 ( .A(ALU_DW01_ash_0__n854), .Y(ALU__N290) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U705 ( .A(ALU_DW01_ash_0__n224), .Y(ALU_DW01_ash_0__n542) );
  O2A1O1Ixp33_ASAP7_75t_R ALU___ALU_DW01_ash_0___U706 ( .A1(ALU_DW01_ash_0__n542), .A2(ALU_DW01_ash_0__n367), .B(ALU_DW01_ash_0__n313), .C(ALU_DW01_ash_0__n551), .Y(
        N289) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U707 ( .A(ALU_DW01_ash_0__n66), .Y(ALU_DW01_ash_0__n699) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U708 ( .A(ALU_DW01_ash_0__n709), .Y(ALU_DW01_ash_0__n698) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U709 ( .A(ALU_DW01_ash_0__n712), .Y(ALU_DW01_ash_0__n697) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U710 ( .A(ALU_DW01_ash_0__n376), .Y(ALU_DW01_ash_0__n708) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U711 ( .A(ALU_DW01_ash_0__n334), .Y(ALU_DW01_ash_0__n696) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U712 ( .A(ALU_DW01_ash_0__n78), .Y(ALU_DW01_ash_0__n720) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U713 ( .A(ALU_DW01_ash_0__n203), .Y(ALU_DW01_ash_0__n719) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U714 ( .A(ALU_DW01_ash_0__n322), .Y(ALU_DW01_ash_0__n718) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U715 ( .A(ALU_DW01_ash_0__n65), .Y(ALU_DW01_ash_0__n717) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U716 ( .A(ALU_DW01_ash_0__n202), .Y(ALU_DW01_ash_0__n721) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U717 ( .A1(ALU_DW01_ash_0__n380), .A2(ALU_DW01_ash_0__n564), .B1(ALU_DW01_ash_0__n612), .B2(ALU_DW01_ash_0__n580), .C(
        n544), .Y(ALU_DW01_ash_0__n772) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U718 ( .A(ALU_DW01_ash_0__n290), .Y(ALU_DW01_ash_0__n543) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U719 ( .A(ALU_DW01_ash_0__n545), .Y(ALU_DW01_ash_0__n544) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U720 ( .A(ALU_DW01_ash_0__n835), .Y(ALU_DW01_ash_0__n545) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U721 ( .A(ALU_DW01_ash_0__n447), .Y(ALU_DW01_ash_0__n546) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U722 ( .A(ALU_DW01_ash_0__n449), .Y(ALU_DW01_ash_0__n547) );
  AND4x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U723 ( .A(ALU_DW01_ash_0__n294), .B(ALU_DW01_ash_0__n484), .C(ALU_DW01_ash_0__n549), .D(ALU_DW01_ash_0__n550), .Y(ALU_DW01_ash_0__n748)
         );
  OR2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U724 ( .A(ALU_DW01_ash_0__n231), .B(ALU_DW01_ash_0__n628), .Y(ALU_DW01_ash_0__n821) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U725 ( .A(n1114), .Y(ALU_DW01_ash_0__n553) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U726 ( .A(n1114), .Y(ALU_DW01_ash_0__n554) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U727 ( .A(n1114), .Y(ALU_DW01_ash_0__n555) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U728 ( .A(ALU_DW01_ash_0__n557), .Y(ALU_DW01_ash_0__n556) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U729 ( .A(ALU_DW01_ash_0__n493), .Y(ALU_DW01_ash_0__n557) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U730 ( .A1(ALU_DW01_ash_0__n663), .A2(n1182), .B1(ALU_DW01_ash_0__n681), .B2(ALU_DW01_ash_0__n536), .C(
        n559), .Y(ALU_DW01_ash_0__n753) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U731 ( .A(ALU_DW01_ash_0__n822), .Y(ALU_DW01_ash_0__n559) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U732 ( .A(ALU_DW01_ash_0__n878), .Y(ALU_DW01_ash_0__n570) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U733 ( .A(ALU_DW01_ash_0__n570), .Y(ALU_DW01_ash_0__n560) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U734 ( .A1(ALU_DW01_ash_0__n522), .A2(ALU_DW01_ash_0__n619), .B1(ALU_DW01_ash_0__n131), .B2(ALU_DW01_ash_0__n331), .C(
        n562), .Y(ALU_DW01_ash_0__n868) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U735 ( .A(ALU_DW01_ash_0__n168), .Y(ALU__N275) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U736 ( .A(ALU_DW01_ash_0__n563), .Y(ALU_DW01_ash_0__n562) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U737 ( .A(ALU_DW01_ash_0__n827), .Y(ALU_DW01_ash_0__n563) );
  AO22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U738 ( .A1(ALU_DW01_ash_0__n688), .A2(n1015), .B1(ALU_DW01_ash_0__n660), .B2(n964), .Y(
        n800) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U739 ( .A1(ALU_DW01_ash_0__n668), .A2(n973), .B1(ALU_DW01_ash_0__n686), .B2(ALU_DW01_ash_0__n554), .C(
        n566), .Y(ALU_DW01_ash_0__n810) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U740 ( .A(ALU_DW01_ash_0__n843), .Y(ALU_DW01_ash_0__n566) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U741 ( .A1(ALU_DW01_ash_0__n664), .A2(ALU_DW01_ash_0__n504), .B1(ALU_DW01_ash_0__n682), .B2(n1182), .C(
        n568), .Y(ALU_DW01_ash_0__n766) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U742 ( .A(ALU_DW01_ash_0__n824), .Y(ALU_DW01_ash_0__n568) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U743 ( .A(ALU_DW01_ash_0__n870), .Y(ALU__N273) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U744 ( .A(ALU_DW01_ash_0__n388), .B(ALU_DW01_ash_0__n621), .Y(ALU_DW01_ash_0__n878) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U745 ( .A(ALU_DW01_ash_0__n201), .Y(ALU_DW01_ash_0__n716) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U746 ( .A(ALU_DW01_ash_0__n204), .Y(ALU_DW01_ash_0__n715) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U747 ( .A(ALU_DW01_ash_0__n321), .Y(ALU_DW01_ash_0__n714) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U748 ( .A(ALU_DW01_ash_0__n43), .Y(ALU_DW01_ash_0__n725) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U749 ( .A1(ALU_DW01_ash_0__n668), .A2(ALU_DW01_ash_0__n555), .B1(ALU_DW01_ash_0__n684), .B2(n929), .C(
        n572), .Y(ALU_DW01_ash_0__n806) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U750 ( .A(ALU_DW01_ash_0__n840), .Y(ALU_DW01_ash_0__n572) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U751 ( .A(ALU_DW01_ash_0__n324), .Y(ALU_DW01_ash_0__n724) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U752 ( .A(ALU_DW01_ash_0__n574), .Y(ALU_DW01_ash_0__n573) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U753 ( .A(ALU_DW01_ash_0__n754), .Y(ALU_DW01_ash_0__n574) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U754 ( .A(n1152), .Y(ALU_DW01_ash_0__n577) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U755 ( .A(n1152), .Y(ALU_DW01_ash_0__n578) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U756 ( .A(n1152), .Y(ALU_DW01_ash_0__n579) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U757 ( .A1(ALU_DW01_ash_0__n667), .A2(ALU_DW01_ash_0__n457), .B1(ALU_DW01_ash_0__n681), .B2(ALU_DW01_ash_0__n259), .C(
        n581), .Y(ALU_DW01_ash_0__n799) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U758 ( .A(ALU_DW01_ash_0__n838), .Y(ALU_DW01_ash_0__n581) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U759 ( .A(ALU_DW01_ash_0__n372), .Y(ALU_DW01_ash_0__n723) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U760 ( .A1(ALU_DW01_ash_0__n660), .A2(n969), .B1(ALU_DW01_ash_0__n678), .B2(n925), .C(
        n583), .Y(ALU_DW01_ash_0__n789) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U761 ( .A(ALU_DW01_ash_0__n241), .Y(ALU_DW01_ash_0__n582) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U762 ( .A(ALU_DW01_ash_0__n832), .Y(ALU_DW01_ash_0__n583) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U763 ( .A1(ALU_DW01_ash_0__n669), .A2(n1029), .B1(ALU_DW01_ash_0__n686), .B2(n1229), .C(
        n585), .Y(ALU_DW01_ash_0__n813) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U764 ( .A(ALU_DW01_ash_0__n844), .Y(ALU_DW01_ash_0__n585) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U765 ( .A(ALU_DW01_ash_0__n376), .Y(ALU_DW01_ash_0__n705) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U766 ( .A(ALU_DW01_ash_0__n777), .Y(ALU_DW01_ash_0__n586) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U767 ( .A(ALU_DW01_ash_0__n376), .Y(ALU_DW01_ash_0__n707) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U768 ( .A(ALU_DW01_ash_0__n733), .Y(ALU_DW01_ash_0__n587) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U769 ( .A(n749), .Y(ALU_DW01_ash_0__n733) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U770 ( .A(ALU_DW01_ash_0__n481), .B(ALU_DW01_ash_0__n621), .Y(ALU_DW01_ash_0__n875) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U771 ( .A(ALU_DW01_ash_0__n343), .B(n749), .Y(ALU_DW01_ash_0__n760) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U772 ( .A(ALU_DW01_ash_0__n631), .B(ALU_DW01_ash_0__n342), .Y(ALU_DW01_ash_0__n757) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U773 ( .A(n964), .B(ALU_DW01_ash_0__n688), .Y(ALU_DW01_ash_0__n805) );
  INVx5_ASAP7_75t_R ALU___ALU_DW01_ash_0___U774 ( .A(ALU_DW01_ash_0__n84), .Y(ALU_DW01_ash_0__n589) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U775 ( .A(ALU_DW01_ash_0__n731), .Y(ALU_DW01_ash_0__n590) );
  OA221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U776 ( .A1(ALU_DW01_ash_0__n380), .A2(ALU_DW01_ash_0__n622), .B1(ALU_DW01_ash_0__n612), .B2(ALU_DW01_ash_0__n603), .C(
        n592), .Y(ALU_DW01_ash_0__n763) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U777 ( .A(ALU_DW01_ash_0__n210), .Y(ALU_DW01_ash_0__n591) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U778 ( .A(ALU_DW01_ash_0__n593), .Y(ALU_DW01_ash_0__n592) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U779 ( .A(ALU_DW01_ash_0__n833), .Y(ALU_DW01_ash_0__n593) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U780 ( .A1(ALU_DW01_ash_0__n664), .A2(n1073), .B1(ALU_DW01_ash_0__n683), .B2(ALU_DW01_ash_0__n504), .C(
        n595), .Y(ALU_DW01_ash_0__n775) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U781 ( .A(ALU_DW01_ash_0__n826), .Y(ALU_DW01_ash_0__n595) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U782 ( .A1(ALU_DW01_ash_0__n661), .A2(n1229), .B1(ALU_DW01_ash_0__n685), .B2(ALU_DW01_ash_0__n578), .C(
        n597), .Y(ALU_DW01_ash_0__n809) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U783 ( .A(ALU_DW01_ash_0__n842), .Y(ALU_DW01_ash_0__n597) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U784 ( .A(ALU_DW01_ash_0__n72), .Y(ALU_DW01_ash_0__n704) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U785 ( .A(ALU_DW01_ash_0__n602), .Y(ALU_DW01_ash_0__n601) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U786 ( .A(ALU_DW01_ash_0__n742), .Y(ALU_DW01_ash_0__n602) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U787 ( .A1(ALU_DW01_ash_0__n665), .A2(ALU_DW01_ash_0__n259), .B1(ALU_DW01_ash_0__n678), .B2(n973), .C(
        n604), .Y(ALU_DW01_ash_0__n814) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U788 ( .A(ALU_DW01_ash_0__n845), .Y(ALU_DW01_ash_0__n604) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U789 ( .A(ALU_DW01_ash_0__n711), .Y(ALU_DW01_ash_0__n701) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U790 ( .A1(ALU_DW01_ash_0__n666), .A2(ALU_DW01_ash_0__n143), .B1(ALU_DW01_ash_0__n678), .B2(n1020), .C(
        n606), .Y(ALU_DW01_ash_0__n798) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U791 ( .A(ALU_DW01_ash_0__n182), .Y(ALU_DW01_ash_0__n605) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U792 ( .A(ALU_DW01_ash_0__n837), .Y(ALU_DW01_ash_0__n606) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U793 ( .A(ALU_DW01_ash_0__n365), .B(ALU_DW01_ash_0__n621), .Y(ALU_DW01_ash_0__n879) );
  AO221x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U794 ( .A1(ALU_DW01_ash_0__n668), .A2(ALU_DW01_ash_0__n579), .B1(ALU_DW01_ash_0__n685), .B2(ALU_DW01_ash_0__n141), .C(
        n610), .Y(ALU_DW01_ash_0__n803) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U795 ( .A(ALU_DW01_ash_0__n841), .Y(ALU_DW01_ash_0__n610) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U796 ( .A(ALU_DW01_ash_0__n207), .Y(ALU_DW01_ash_0__n703) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U797 ( .A(ALU_DW01_ash_0__n345), .Y(ALU_DW01_ash_0__n611) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U798 ( .A(ALU_DW01_ash_0__n385), .Y(ALU_DW01_ash_0__n612) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U799 ( .A(ALU_DW01_ash_0__n387), .Y(ALU_DW01_ash_0__n613) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U800 ( .A(ALU_DW01_ash_0__n735), .B(ALU_DW01_ash_0__n508), .Y(ALU_DW01_ash_0__n752) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U801 ( .A(ALU_DW01_ash_0__n575), .B(ALU_DW01_ash_0__n621), .Y(ALU_DW01_ash_0__n876) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U802 ( .A(ALU_DW01_ash_0__n369), .Y(ALU_DW01_ash_0__n673) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U803 ( .A(ALU_DW01_ash_0__n615), .Y(ALU_DW01_ash_0__n680) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U804 ( .A(ALU_DW01_ash_0__n690), .Y(ALU_DW01_ash_0__n678) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U805 ( .A(ALU_DW01_ash_0__n734), .B(ALU_DW01_ash_0__n735), .Y(ALU_DW01_ash_0__n617) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U806 ( .A(ALU_DW01_ash_0__n573), .Y(ALU_DW01_ash_0__n618) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U807 ( .A(ALU_DW01_ash_0__n507), .Y(ALU_DW01_ash_0__n734) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U808 ( .A(ALU_DW01_ash_0__n450), .B(ALU_DW01_ash_0__n508), .Y(ALU_DW01_ash_0__n790) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U809 ( .A(ALU_DW01_ash_0__n599), .B(ALU_DW01_ash_0__n621), .Y(ALU_DW01_ash_0__n877) );
  AO222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U810 ( .A1(ALU_DW01_ash_0__n660), .A2(n1015), .B1(n964), .B2(ALU_DW01_ash_0__n696), .C1(
        n686), .C2(ALU_DW01_ash_0__n427), .Y(ALU_DW01_ash_0__n769) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U811 ( .A(ALU_DW01_ash_0__n671), .Y(ALU_DW01_ash_0__n670) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U812 ( .A(ALU_DW01_ash_0__n671), .Y(ALU_DW01_ash_0__n669) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U813 ( .A(ALU_DW01_ash_0__n28), .Y(ALU_DW01_ash_0__n671) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U814 ( .A(ALU_DW01_ash_0__n318), .Y(ALU_DW01_ash_0__n675) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U815 ( .A(ALU_DW01_ash_0__n677), .Y(ALU_DW01_ash_0__n676) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U816 ( .A(ALU_DW01_ash_0__n60), .Y(ALU_DW01_ash_0__n695) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U817 ( .A(ALU_DW01_ash_0__n451), .B(ALU_DW01_ash_0__n734), .Y(ALU_DW01_ash_0__n792) );
  AND2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U818 ( .A(ALU_DW01_ash_0__n735), .B(ALU_DW01_ash_0__n508), .Y(ALU_DW01_ash_0__n756) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U819 ( .A(ALU_DW01_ash_0__n408), .Y(ALU_DW01_ash_0__n736) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_ash_0___U820 ( .A(ALU_DW01_ash_0__n71), .Y(ALU_DW01_ash_0__n626) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U821 ( .A(ALU_DW01_ash_0__n173), .Y(ALU_DW01_ash_0__n627) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U822 ( .A(ALU_DW01_ash_0__n304), .Y(ALU_DW01_ash_0__n628) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U823 ( .A(ALU_DW01_ash_0__n410), .B(ALU_DW01_ash_0__n628), .Y(ALU_DW01_ash_0__n746) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U824 ( .A(ALU_DW01_ash_0__n335), .B(ALU_DW01_ash_0__n621), .Y(ALU_DW01_ash_0__n872) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U825 ( .A(ALU_DW01_ash_0__n589), .B(ALU_DW01_ash_0__n332), .Y(ALU_DW01_ash_0__n884) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U826 ( .A(ALU_DW01_ash_0__n524), .Y(ALU__N259) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U827 ( .A(ALU_DW01_ash_0__n638), .Y(ALU_DW01_ash_0__n635) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U828 ( .A(ALU_DW01_ash_0__n54), .Y(ALU_DW01_ash_0__n636) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_ash_0___U829 ( .A(ALU_DW01_ash_0__n639), .Y(ALU_DW01_ash_0__n638) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_ash_0___U830 ( .A(ALU_DW01_ash_0__n351), .Y(ALU_DW01_ash_0__n639) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U831 ( .A(ALU_DW01_ash_0__n208), .Y(ALU_DW01_ash_0__n700) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U832 ( .A(ALU_DW01_ash_0__n123), .Y(ALU_DW01_ash_0__n643) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U833 ( .A(ALU_DW01_ash_0__n153), .Y(ALU_DW01_ash_0__n650) );
  OR2x6_ASAP7_75t_R ALU___ALU_DW01_ash_0___U834 ( .A(ALU_DW01_ash_0__n621), .B(ALU_DW01_ash_0__n628), .Y(ALU_DW01_ash_0__n744) );
  O2A1O1Ixp33_ASAP7_75t_R ALU___ALU_DW01_ash_0___U835 ( .A1(ALU_DW01_ash_0__n500), .A2(ALU_DW01_ash_0__n367), .B(ALU_DW01_ash_0__n421), .C(ALU_DW01_ash_0__n551), .Y(
        n854) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U836 ( .A1(ALU_DW01_ash_0__n708), .A2(n1215), .B1(ALU_DW01_ash_0__n725), .B2(n920), .Y(
        n758) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U837 ( .A1(ALU_DW01_ash_0__n707), .A2(n920), .B1(ALU_DW01_ash_0__n714), .B2(n1160), .Y(
        n768) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U838 ( .A1(ALU_DW01_ash_0__n707), .A2(n1160), .B1(ALU_DW01_ash_0__n714), .B2(n1100), .Y(
        n777) );
  O2A1O1Ixp33_ASAP7_75t_R ALU___ALU_DW01_ash_0___U839 ( .A1(ALU_DW01_ash_0__n456), .A2(ALU_DW01_ash_0__n367), .B(ALU_DW01_ash_0__n513), .C(ALU_DW01_ash_0__n551), .Y(
        n856) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U840 ( .A1(ALU_DW01_ash_0__n626), .A2(ALU_DW01_ash_0__n335), .B1(ALU_DW01_ash_0__n85), .B2(ALU_DW01_ash_0__n233), .Y(ALU_DW01_ash_0__n779) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U841 ( .A1(ALU_DW01_ash_0__n491), .A2(ALU_DW01_ash_0__n611), .B1(ALU_DW01_ash_0__n131), .B2(ALU_DW01_ash_0__n380), .C1(
        n444), .C2(ALU_DW01_ash_0__n461), .Y(ALU_DW01_ash_0__n781) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U842 ( .A1(ALU_DW01_ash_0__n582), .A2(ALU_DW01_ash_0__n619), .B1(ALU_DW01_ash_0__n477), .B2(ALU_DW01_ash_0__n539), .C1(
        n558), .C2(ALU_DW01_ash_0__n196), .Y(ALU_DW01_ash_0__n788) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U843 ( .A1(ALU_DW01_ash_0__n114), .A2(ALU_DW01_ash_0__n619), .B1(ALU_DW01_ash_0__n520), .B2(ALU_DW01_ash_0__n539), .C1(
        n567), .C2(ALU_DW01_ash_0__n197), .Y(ALU_DW01_ash_0__n795) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U844 ( .A1(ALU_DW01_ash_0__n605), .A2(ALU_DW01_ash_0__n619), .B1(ALU_DW01_ash_0__n509), .B2(ALU_DW01_ash_0__n539), .C1(
        n594), .C2(ALU_DW01_ash_0__n196), .Y(ALU_DW01_ash_0__n797) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U845 ( .A1(ALU_DW01_ash_0__n580), .A2(ALU_DW01_ash_0__n460), .B1(ALU_DW01_ash_0__n564), .B2(ALU_DW01_ash_0__n612), .C1(
        n145), .C2(ALU_DW01_ash_0__n627), .Y(ALU_DW01_ash_0__n737) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U846 ( .A1(n1024), .A2(ALU_DW01_ash_0__n722), .B1(ALU_DW01_ash_0__n503), .B2(ALU_DW01_ash_0__n697), .Y(
        n801) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U847 ( .A1(ALU_DW01_ash_0__n609), .A2(ALU_DW01_ash_0__n619), .B1(ALU_DW01_ash_0__n491), .B2(ALU_DW01_ash_0__n539), .C1(
        n131), .C2(ALU_DW01_ash_0__n197), .Y(ALU_DW01_ash_0__n802) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U848 ( .A1(ALU_DW01_ash_0__n522), .A2(ALU_DW01_ash_0__n460), .B1(ALU_DW01_ash_0__n611), .B2(ALU_DW01_ash_0__n589), .C1(
        n571), .C2(ALU_DW01_ash_0__n627), .Y(ALU_DW01_ash_0__n738) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U849 ( .A1(ALU_DW01_ash_0__n189), .A2(ALU_DW01_ash_0__n725), .B1(n1024), .B2(ALU_DW01_ash_0__n697), .Y(
        n807) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U850 ( .A1(ALU_DW01_ash_0__n596), .A2(ALU_DW01_ash_0__n619), .B1(ALU_DW01_ash_0__n558), .B2(ALU_DW01_ash_0__n539), .C1(
        n582), .C2(ALU_DW01_ash_0__n197), .Y(ALU_DW01_ash_0__n808) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U851 ( .A1(ALU_DW01_ash_0__n565), .A2(ALU_DW01_ash_0__n552), .B1(ALU_DW01_ash_0__n401), .B2(ALU_DW01_ash_0__n460), .Y(
        n739) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U852 ( .A1(n1068), .A2(ALU_DW01_ash_0__n717), .B1(ALU_DW01_ash_0__n192), .B2(ALU_DW01_ash_0__n698), .Y(
        n811) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U853 ( .A1(ALU_DW01_ash_0__n584), .A2(ALU_DW01_ash_0__n301), .B1(ALU_DW01_ash_0__n567), .B2(ALU_DW01_ash_0__n538), .C1(
        n115), .C2(ALU_DW01_ash_0__n197), .Y(ALU_DW01_ash_0__n812) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U854 ( .A1(ALU_DW01_ash_0__n603), .A2(ALU_DW01_ash_0__n552), .B1(ALU_DW01_ash_0__n622), .B2(ALU_DW01_ash_0__n462), .Y(
        n740) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U855 ( .A1(ALU_DW01_ash_0__n144), .A2(ALU_DW01_ash_0__n619), .B1(ALU_DW01_ash_0__n594), .B2(ALU_DW01_ash_0__n538), .C1(
        n605), .C2(ALU_DW01_ash_0__n197), .Y(ALU_DW01_ash_0__n816) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U856 ( .A1(ALU_DW01_ash_0__n580), .A2(ALU_DW01_ash_0__n627), .B1(ALU_DW01_ash_0__n564), .B2(ALU_DW01_ash_0__n462), .Y(
        n741) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U857 ( .A1(ALU_DW01_ash_0__n504), .A2(ALU_DW01_ash_0__n718), .B1(n1182), .B2(ALU_DW01_ash_0__n699), .Y(
        n819) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U858 ( .A1(ALU_DW01_ash_0__n196), .A2(ALU_DW01_ash_0__n596), .B1(ALU_DW01_ash_0__n212), .B2(ALU_DW01_ash_0__n401), .C1(
        n538), .C2(ALU_DW01_ash_0__n582), .Y(ALU_DW01_ash_0__n820) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U859 ( .A1(n1073), .A2(ALU_DW01_ash_0__n719), .B1(ALU_DW01_ash_0__n504), .B2(ALU_DW01_ash_0__n696), .Y(
        n822) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U860 ( .A1(ALU_DW01_ash_0__n196), .A2(ALU_DW01_ash_0__n584), .B1(ALU_DW01_ash_0__n212), .B2(ALU_DW01_ash_0__n622), .C1(
        n538), .C2(ALU_DW01_ash_0__n115), .Y(ALU_DW01_ash_0__n823) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U861 ( .A1(n925), .A2(ALU_DW01_ash_0__n720), .B1(n1073), .B2(ALU_DW01_ash_0__n708), .Y(
        n824) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U862 ( .A1(ALU_DW01_ash_0__n196), .A2(ALU_DW01_ash_0__n144), .B1(ALU_DW01_ash_0__n212), .B2(ALU_DW01_ash_0__n564), .C1(
        n538), .C2(ALU_DW01_ash_0__n605), .Y(ALU_DW01_ash_0__n825) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U863 ( .A1(n969), .A2(ALU_DW01_ash_0__n720), .B1(n925), .B2(ALU_DW01_ash_0__n700), .Y(
        n826) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U864 ( .A1(ALU_DW01_ash_0__n196), .A2(ALU_DW01_ash_0__n571), .B1(ALU_DW01_ash_0__n212), .B2(ALU_DW01_ash_0__n589), .C1(
        n538), .C2(ALU_DW01_ash_0__n609), .Y(ALU_DW01_ash_0__n827) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U865 ( .A1(ALU_DW01_ash_0__n47), .A2(ALU_DW01_ash_0__n721), .B1(n969), .B2(ALU_DW01_ash_0__n700), .Y(
        n829) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U866 ( .A(ALU_DW01_ash_0__n517), .B(ALU_DW01_ash_0__n607), .Y(ALU_DW01_ash_0__n869) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U867 ( .A1(ALU_DW01_ash_0__n582), .A2(ALU_DW01_ash_0__n552), .B1(ALU_DW01_ash_0__n596), .B2(ALU_DW01_ash_0__n461), .Y(
        n831) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U868 ( .A(ALU_DW01_ash_0__n591), .B(ALU_DW01_ash_0__n607), .Y(ALU_DW01_ash_0__n870) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U869 ( .A1(ALU_DW01_ash_0__n114), .A2(ALU_DW01_ash_0__n552), .B1(ALU_DW01_ash_0__n584), .B2(ALU_DW01_ash_0__n461), .Y(
        n833) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U870 ( .A(ALU_DW01_ash_0__n543), .B(ALU_DW01_ash_0__n607), .Y(ALU_DW01_ash_0__n871) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U871 ( .A1(ALU_DW01_ash_0__n605), .A2(ALU_DW01_ash_0__n627), .B1(ALU_DW01_ash_0__n145), .B2(ALU_DW01_ash_0__n462), .Y(
        n835) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U872 ( .A1(n1229), .A2(ALU_DW01_ash_0__n723), .B1(ALU_DW01_ash_0__n578), .B2(ALU_DW01_ash_0__n333), .Y(
        n837) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U873 ( .A(ALU_DW01_ash_0__n734), .B(ALU_DW01_ash_0__n735), .Y(ALU_DW01_ash_0__n754) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U874 ( .A1(ALU_DW01_ash_0__n627), .A2(ALU_DW01_ash_0__n609), .B1(ALU_DW01_ash_0__n461), .B2(ALU_DW01_ash_0__n571), .C1(
        n735), .C2(ALU_DW01_ash_0__n601), .Y(ALU_DW01_ash_0__n780) );
  OA22x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U875 ( .A1(ALU_DW01_ash_0__n508), .A2(ALU_DW01_ash_0__n522), .B1(ALU_DW01_ash_0__n734), .B2(ALU_DW01_ash_0__n589), .Y(
        n742) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U876 ( .A1(ALU_DW01_ash_0__n259), .A2(ALU_DW01_ash_0__n724), .B1(n973), .B2(ALU_DW01_ash_0__n703), .Y(
        n840) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U877 ( .A1(n1029), .A2(ALU_DW01_ash_0__n724), .B1(n1229), .B2(ALU_DW01_ash_0__n703), .Y(
        n841) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U878 ( .A1(ALU_DW01_ash_0__n565), .A2(ALU_DW01_ash_0__n460), .B1(ALU_DW01_ash_0__n401), .B2(ALU_DW01_ash_0__n612), .C1(
        n596), .C2(ALU_DW01_ash_0__n552), .Y(ALU_DW01_ash_0__n786) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U879 ( .A1(n929), .A2(ALU_DW01_ash_0__n725), .B1(n1029), .B2(ALU_DW01_ash_0__n704), .Y(
        n842) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U880 ( .A1(ALU_DW01_ash_0__n457), .A2(ALU_DW01_ash_0__n725), .B1(ALU_DW01_ash_0__n259), .B2(ALU_DW01_ash_0__n704), .Y(
        n843) );
  OA222x2_ASAP7_75t_R ALU___ALU_DW01_ash_0___U881 ( .A1(ALU_DW01_ash_0__n603), .A2(ALU_DW01_ash_0__n460), .B1(ALU_DW01_ash_0__n622), .B2(ALU_DW01_ash_0__n612), .C1(
        n584), .C2(ALU_DW01_ash_0__n254), .Y(ALU_DW01_ash_0__n794) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U882 ( .A1(ALU_DW01_ash_0__n554), .A2(ALU_DW01_ash_0__n715), .B1(n929), .B2(ALU_DW01_ash_0__n705), .Y(
        n844) );
  AO22x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U883 ( .A1(n1060), .A2(ALU_DW01_ash_0__n719), .B1(ALU_DW01_ash_0__n457), .B2(ALU_DW01_ash_0__n701), .Y(
        n845) );
  OR3x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U884 ( .A(n798), .B(n888), .C(ALU_DW01_ash_0__n364), .Y(ALU_DW01_ash_0__n850) );
  OR3x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U885 ( .A(n851), .B(n955), .C(n1056), .Y(ALU_DW01_ash_0__n851) );
  OR3x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U886 ( .A(ALU_DW01_ash_0__n319), .B(n790), .C(n547), .Y(ALU_DW01_ash_0__n852) );
  OR3x1_ASAP7_75t_R ALU___ALU_DW01_ash_0___U887 ( .A(n1222), .B(n794), .C(n767), .Y(ALU_DW01_ash_0__n853) );

  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_31 ( .A(ALU_DW01_sub_0__n697), .B(n1091), .CI(ALU_DW01_sub_0__n637), .SN(ALU_DW01_sub_0__n705) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_29 ( .A(n1215), .B(ALU_DW01_sub_0__n614), .CI(ALU_DW01_sub_0__n613), .CON(ALU_DW01_sub_0__n706), .SN(
        n707) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_28 ( .A(n920), .B(ALU_DW01_sub_0__n525), .CI(ALU_DW01_sub_0__n649), .CON(ALU_DW01_sub_0__n708), .SN(
        n709) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_27 ( .A(ALU_DW01_sub_0__n645), .B(n1160), .CI(ALU_DW01_sub_0__n644), .CON(ALU_DW01_sub_0__n710), .SN(
        n711) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_26 ( .A(n1100), .B(ALU_DW01_sub_0__n378), .CI(ALU_DW01_sub_0__n651), .CON(ALU_DW01_sub_0__n712), .SN(
        n713) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_24 ( .A(n1064), .B(ALU_DW01_sub_0__n600), .CI(ALU_DW01_sub_0__n599), .CON(ALU_DW01_sub_0__n714), .SN(
        n715) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_22 ( .A(n1024), .B(ALU_DW01_sub_0__n563), .CI(ALU_DW01_sub_0__n655), .CON(ALU_DW01_sub_0__n716), .SN(
        n717) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_21 ( .A(ALU_DW01_sub_0__n588), .B(n1225), .CI(ALU_DW01_sub_0__n587), .CON(ALU_DW01_sub_0__n718), .SN(
        n719) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_20 ( .A(n1068), .B(ALU_DW01_sub_0__n575), .CI(ALU_DW01_sub_0__n574), .CON(ALU_DW01_sub_0__n720), .SN(
        n721) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_18 ( .A(ALU_DW01_sub_0__n617), .B(ALU_DW01_sub_0__n618), .CI(n1182), .CON(ALU_DW01_sub_0__n722), .SN(
        n723) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_16 ( .A(ALU_DW01_sub_0__n680), .B(n1073), .CI(ALU_DW01_sub_0__n660), .CON(ALU_DW01_sub_0__n724), .SN(
        n725) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_15 ( .A(n925), .B(ALU_DW01_sub_0__n604), .CI(ALU_DW01_sub_0__n603), .CON(ALU_DW01_sub_0__n726), .SN(
        n727) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_14 ( .A(ALU_DW01_sub_0__n296), .B(n969), .CI(ALU_DW01_sub_0__n661), .CON(ALU_DW01_sub_0__n728), .SN(
        n729) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_13 ( .A(n1020), .B(ALU_DW01_sub_0__n677), .CI(ALU_DW01_sub_0__n621), .CON(ALU_DW01_sub_0__n730), .SN(
        n731) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_12 ( .A(ALU_DW01_sub_0__n676), .B(n1109), .CI(ALU_DW01_sub_0__n662), .CON(ALU_DW01_sub_0__n732), .SN(
        n733) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_11 ( .A(ALU_DW01_sub_0__n663), .B(ALU_DW01_sub_0__n607), .CI(n1152), .CON(ALU_DW01_sub_0__n734), .SN(
        n735) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_10 ( .A(ALU_DW01_sub_0__n624), .B(n1229), .CI(ALU_DW01_sub_0__n664), .CON(ALU_DW01_sub_0__n736), .SN(
        n737) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_9 ( .A(ALU_DW01_sub_0__n632), .B(n1029), .CI(ALU_DW01_sub_0__n631), .CON(ALU_DW01_sub_0__n738), .SN(ALU_DW01_sub_0__n739)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_8 ( .A(n929), .B(ALU_DW01_sub_0__n450), .CI(ALU_DW01_sub_0__n666), .CON(ALU_DW01_sub_0__n740), .SN(ALU_DW01_sub_0__n741)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_7 ( .A(ALU_DW01_sub_0__n635), .B(ALU_DW01_sub_0__n636), .CI(n1114), .CON(ALU_DW01_sub_0__n742), .SN(ALU_DW01_sub_0__n743)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_6 ( .A(n973), .B(ALU_DW01_sub_0__n609), .CI(ALU_DW01_sub_0__n668), .CON(ALU_DW01_sub_0__n744), .SN(ALU_DW01_sub_0__n745)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_5 ( .A(ALU_DW01_sub_0__n628), .B(n1233), .CI(ALU_DW01_sub_0__n627), .CON(ALU_DW01_sub_0__n746), .SN(ALU_DW01_sub_0__n747)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_3 ( .A(n1060), .B(ALU_DW01_sub_0__n592), .CI(ALU_DW01_sub_0__n591), .CON(ALU_DW01_sub_0__n748), .SN(ALU_DW01_sub_0__n749)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2_1 ( .A(n1015), .B(ALU_DW01_sub_0__n579), .CI(ALU_DW01_sub_0__n521), .CON(ALU_DW01_sub_0__n750), .SN(ALU_DW01_sub_0__n751)
         );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U1 ( .A(ALU_DW01_sub_0__n737), .Y(ALU_DW01_sub_0__n1) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U2 ( .A(ALU_DW01_sub_0__n731), .Y(ALU_DW01_sub_0__n2) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U3 ( .A(ALU_DW01_sub_0__n729), .Y(ALU_DW01_sub_0__n3) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U4 ( .A(ALU_DW01_sub_0__n727), .Y(ALU_DW01_sub_0__n4) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U5 ( .A(ALU_DW01_sub_0__n707), .Y(ALU_DW01_sub_0__n5) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U6 ( .A(ALU_DW01_sub_0__n751), .Y(ALU_DW01_sub_0__n6) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U7 ( .A(ALU_DW01_sub_0__ALU_DW01_sub_0__n735), .Y(ALU_DW01_sub_0__n7) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U8 ( .A(ALU_DW01_sub_0__n742), .Y(ALU_DW01_sub_0__n8) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_sub_0___U9 ( .A(ALU_DW01_sub_0__n332), .Y(ALU_DW01_sub_0__n635) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U10 ( .A(ALU_DW01_sub_0__n718), .Y(ALU_DW01_sub_0__n9) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U11 ( .A(ALU_DW01_sub_0__n746), .Y(ALU_DW01_sub_0__n10) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U12 ( .A(ALU_DW01_sub_0__n736), .Y(ALU_DW01_sub_0__n11) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U13 ( .A(ALU_DW01_sub_0__n728), .Y(ALU_DW01_sub_0__n12) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U14 ( .A(ALU_DW01_sub_0__n710), .Y(ALU_DW01_sub_0__n13) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U15 ( .A(ALU_DW01_sub_0__n738), .Y(ALU_DW01_sub_0__n14) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U16 ( .A(ALU_DW01_sub_0__n734), .Y(ALU_DW01_sub_0__n15) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U17 ( .A(ALU_DW01_sub_0__n750), .Y(ALU_DW01_sub_0__n16) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U18 ( .A(ALU_DW01_sub_0__n724), .Y(ALU_DW01_sub_0__n17) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U19 ( .A(ALU_DW01_sub_0__n732), .Y(ALU_DW01_sub_0__n18) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U20 ( .A(ALU_DW01_sub_0__n730), .Y(ALU_DW01_sub_0__n19) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U21 ( .A(ALU_DW01_sub_0__n726), .Y(ALU_DW01_sub_0__n20) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U22 ( .A(ALU_DW01_sub_0__n740), .Y(ALU_DW01_sub_0__n21) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U23 ( .A(ALU_DW01_sub_0__n716), .Y(ALU_DW01_sub_0__n22) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U24 ( .A(ALU_DW01_sub_0__n714), .Y(ALU_DW01_sub_0__n23) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U25 ( .A(ALU_DW01_sub_0__n744), .Y(ALU_DW01_sub_0__n24) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U26 ( .A(ALU_DW01_sub_0__n708), .Y(ALU_DW01_sub_0__n25) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U27 ( .A(ALU_DW01_sub_0__n748), .Y(ALU_DW01_sub_0__n26) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U28 ( .A(ALU_DW01_sub_0__n712), .Y(ALU_DW01_sub_0__n27) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U29 ( .A(ALU_DW01_sub_0__n720), .Y(ALU_DW01_sub_0__n28) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U30 ( .A(ALU_DW01_sub_0__n706), .Y(ALU_DW01_sub_0__n29) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U31 ( .A(ALU_DW01_sub_0__n722), .Y(ALU_DW01_sub_0__n30) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U32 ( .A(ALU_DW01_sub_0__n594), .Y(ALU_DW01_sub_0__n617) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U33 ( .A(ALU_DW01_sub_0__n121), .Y(ALU__N176) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U34 ( .A(ALU_DW01_sub_0__n43), .Y(ALU__N169) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U35 ( .A(ALU_DW01_sub_0__n36), .Y(ALU_DW01_sub_0__n121) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U36 ( .A(ALU_DW01_sub_0__n756), .Y(ALU_DW01_sub_0__n33) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U37 ( .A(ALU_DW01_sub_0__n35), .Y(ALU__N177) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U38 ( .A(ALU_DW01_sub_0__n33), .Y(ALU_DW01_sub_0__n35) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U39 ( .A(ALU_DW01_sub_0__n236), .Y(ALU__N174) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U40 ( .A(ALU_DW01_sub_0__n37), .Y(ALU_DW01_sub_0__n236) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U41 ( .A(ALU_DW01_sub_0__n757), .Y(ALU_DW01_sub_0__n36) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U42 ( .A(ALU_DW01_sub_0__n759), .Y(ALU_DW01_sub_0__n37) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U43 ( .A(ALU_DW01_sub_0__n762), .Y(ALU_DW01_sub_0__n38) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U44 ( .A(ALU_DW01_sub_0__n42), .Y(ALU__N171) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U45 ( .A(ALU_DW01_sub_0__n38), .Y(ALU_DW01_sub_0__n42) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U46 ( .A(ALU_DW01_sub_0__n87), .Y(ALU__N173) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U47 ( .A(ALU_DW01_sub_0__n78), .Y(ALU__N175) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U48 ( .A(ALU_DW01_sub_0__n761), .Y(ALU_DW01_sub_0__n41) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U49 ( .A(ALU_DW01_sub_0__n97), .Y(ALU__N159) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U50 ( .A(ALU_DW01_sub_0__n190), .Y(ALU_DW01_sub_0__n764) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U51 ( .A(ALU_DW01_sub_0__n764), .Y(ALU_DW01_sub_0__n43) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U52 ( .A(ALU_DW01_sub_0__n765), .Y(ALU_DW01_sub_0__n44) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U53 ( .A(ALU_DW01_sub_0__n771), .Y(ALU_DW01_sub_0__n45) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U54 ( .A(ALU_DW01_sub_0__n63), .Y(ALU__N162) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U55 ( .A(ALU_DW01_sub_0__n45), .Y(ALU_DW01_sub_0__n63) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U56 ( .A(ALU_DW01_sub_0__n65), .Y(ALU__N170) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U57 ( .A(ALU_DW01_sub_0__n100), .Y(ALU__N167) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U58 ( .A(ALU__n73), .Y(ALU_DW01_sub_0__n701) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U59 ( .A(ALU_DW01_sub_0__ALU_DW01_sub_0__n470), .Y(ALU_DW01_sub_0__n47) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U60 ( .A(ALU_DW01_sub_0__n458), .Y(ALU_DW01_sub_0__n48) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U61 ( .A(ALU_DW01_sub_0__n460), .Y(ALU_DW01_sub_0__n49) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U62 ( .A(ALU_DW01_sub_0__n467), .Y(ALU_DW01_sub_0__n50) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U63 ( .A(ALU_DW01_sub_0__n471), .Y(ALU_DW01_sub_0__n51) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U64 ( .A(ALU_DW01_sub_0__n461), .Y(ALU_DW01_sub_0__n52) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U65 ( .A(ALU_DW01_sub_0__n463), .Y(ALU_DW01_sub_0__n53) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U66 ( .A(ALU_DW01_sub_0__n472), .Y(ALU_DW01_sub_0__n455) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U67 ( .A(ALU_DW01_sub_0__n767), .Y(ALU_DW01_sub_0__n54) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U68 ( .A(ALU_DW01_sub_0__n775), .Y(ALU_DW01_sub_0__n55) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U69 ( .A(ALU_DW01_sub_0__n134), .Y(ALU__N158) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U70 ( .A(ALU_DW01_sub_0__n55), .Y(ALU_DW01_sub_0__n134) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U71 ( .A(ALU_DW01_sub_0__n776), .Y(ALU_DW01_sub_0__n56) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U72 ( .A(ALU_DW01_sub_0__n167), .Y(ALU__N157) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U73 ( .A(ALU_DW01_sub_0__n56), .Y(ALU_DW01_sub_0__n167) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U74 ( .A(ALU_DW01_sub_0__n335), .Y(ALU__N180) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U75 ( .A(ALU_DW01_sub_0__n374), .Y(ALU_DW01_sub_0__n57) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U76 ( .A(ALU_DW01_sub_0__n361), .Y(ALU_DW01_sub_0__n58) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U77 ( .A(ALU_DW01_sub_0__n363), .Y(ALU_DW01_sub_0__n59) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U78 ( .A(ALU_DW01_sub_0__n375), .Y(ALU_DW01_sub_0__n60) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U79 ( .A(ALU_DW01_sub_0__n365), .Y(ALU_DW01_sub_0__n61) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U80 ( .A(ALU_DW01_sub_0__n367), .Y(ALU_DW01_sub_0__n62) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U81 ( .A(ALU_DW01_sub_0__n348), .Y(ALU__N181) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U82 ( .A(ALU_DW01_sub_0__n763), .Y(ALU_DW01_sub_0__n65) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U83 ( .A(ALU_DW01_sub_0__n328), .Y(ALU_DW01_sub_0__n66) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U84 ( .A(ALU_DW01_sub_0__n315), .Y(ALU_DW01_sub_0__n67) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U85 ( .A(ALU_DW01_sub_0__n317), .Y(ALU_DW01_sub_0__n68) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U86 ( .A(ALU_DW01_sub_0__n329), .Y(ALU_DW01_sub_0__n69) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U87 ( .A(ALU_DW01_sub_0__n319), .Y(ALU_DW01_sub_0__n70) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U88 ( .A(ALU_DW01_sub_0__n321), .Y(ALU_DW01_sub_0__n71) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U89 ( .A(ALU_DW01_sub_0__n659), .Y(ALU_DW01_sub_0__n313) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U90 ( .A(ALU_DW01_sub_0__n777), .Y(ALU_DW01_sub_0__n72) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U91 ( .A(ALU_DW01_sub_0__n448), .Y(ALU__N156) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U92 ( .A(ALU_DW01_sub_0__n72), .Y(ALU_DW01_sub_0__n448) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U93 ( .A(ALU_DW01_sub_0__n128), .Y(ALU__N154) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U94 ( .A(ALU_DW01_sub_0__n75), .Y(ALU_DW01_sub_0__n74) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U95 ( .A(ALU_DW01_sub_0__n781), .Y(ALU_DW01_sub_0__n75) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U96 ( .A(ALU_DW01_sub_0__n77), .Y(ALU_DW01_sub_0__n76) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U97 ( .A(ALU_DW01_sub_0__n754), .Y(ALU_DW01_sub_0__n77) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U98 ( .A(ALU_DW01_sub_0__n753), .Y(ALU_DW01_sub_0__n348) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U99 ( .A(ALU_DW01_sub_0__n175), .Y(ALU_DW01_sub_0__n758) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U100 ( .A(ALU_DW01_sub_0__n758), .Y(ALU_DW01_sub_0__n78) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U101 ( .A(ALU_DW01_sub_0__n778), .Y(ALU_DW01_sub_0__n79) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U102 ( .A(ALU_DW01_sub_0__n120), .Y(ALU__N155) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U103 ( .A(ALU_DW01_sub_0__n79), .Y(ALU_DW01_sub_0__n120) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U104 ( .A(ALU_DW01_sub_0__n425), .Y(ALU_DW01_sub_0__n80) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U105 ( .A(ALU_DW01_sub_0__n412), .Y(ALU_DW01_sub_0__n81) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U106 ( .A(ALU_DW01_sub_0__n414), .Y(ALU_DW01_sub_0__n82) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U107 ( .A(ALU_DW01_sub_0__n426), .Y(ALU_DW01_sub_0__n83) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U108 ( .A(ALU_DW01_sub_0__n416), .Y(ALU_DW01_sub_0__n84) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U109 ( .A(ALU_DW01_sub_0__n418), .Y(ALU_DW01_sub_0__n85) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U110 ( .A(ALU_DW01_sub_0__n658), .Y(ALU_DW01_sub_0__n410) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U111 ( .A(ALU_DW01_sub_0__n705), .Y(ALU_DW01_sub_0__n86) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U112 ( .A(ALU_DW01_sub_0__n349), .Y(ALU_DW01_sub_0__n753) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U113 ( .A(ALU_DW01_sub_0__n297), .Y(ALU_DW01_sub_0__n760) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U114 ( .A(ALU_DW01_sub_0__n760), .Y(ALU_DW01_sub_0__n87) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U115 ( .A(ALU_DW01_sub_0__n377), .Y(ALU_DW01_sub_0__n88) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U116 ( .A(ALU_DW01_sub_0__n90), .Y(ALU_DW01_sub_0__n89) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U117 ( .A(ALU_DW01_sub_0__n218), .Y(ALU_DW01_sub_0__n90) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U118 ( .A(ALU_DW01_sub_0__n495), .Y(ALU_DW01_sub_0__n91) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U119 ( .A(ALU_DW01_sub_0__n482), .Y(ALU_DW01_sub_0__n92) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U120 ( .A(ALU_DW01_sub_0__n484), .Y(ALU_DW01_sub_0__n93) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U121 ( .A(ALU_DW01_sub_0__n496), .Y(ALU_DW01_sub_0__n94) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U122 ( .A(ALU_DW01_sub_0__n486), .Y(ALU_DW01_sub_0__n95) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U123 ( .A(ALU_DW01_sub_0__n488), .Y(ALU_DW01_sub_0__n96) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U124 ( .A(ALU_DW01_sub_0__n672), .Y(ALU_DW01_sub_0__n480) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U125 ( .A(ALU_DW01_sub_0__n774), .Y(ALU_DW01_sub_0__n97) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U126 ( .A(ALU_DW01_sub_0__n780), .Y(ALU_DW01_sub_0__n98) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U127 ( .A(ALU_DW01_sub_0__n5), .Y(ALU_DW01_sub_0__n754) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U128 ( .A(ALU_DW01_sub_0__n76), .Y(ALU__N179) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U129 ( .A(ALU_DW01_sub_0__n227), .Y(ALU_DW01_sub_0__n766) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U130 ( .A(ALU_DW01_sub_0__n766), .Y(ALU_DW01_sub_0__n100) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U131 ( .A(ALU_DW01_sub_0__n452), .Y(ALU_DW01_sub_0__n101) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U132 ( .A(ALU_DW01_sub_0__n453), .Y(ALU_DW01_sub_0__n102) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U133 ( .A(ALU_DW01_sub_0__n465), .Y(ALU_DW01_sub_0__n103) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U134 ( .A(ALU_DW01_sub_0__n478), .Y(ALU_DW01_sub_0__n104) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U135 ( .A(ALU_DW01_sub_0__n490), .Y(ALU_DW01_sub_0__n105) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U136 ( .A(ALU_DW01_sub_0__n555), .Y(ALU_DW01_sub_0__n106) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U137 ( .A(ALU_DW01_sub_0__n542), .Y(ALU_DW01_sub_0__n107) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U138 ( .A(ALU_DW01_sub_0__n544), .Y(ALU_DW01_sub_0__n108) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U139 ( .A(ALU_DW01_sub_0__n556), .Y(ALU_DW01_sub_0__n109) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U140 ( .A(ALU_DW01_sub_0__n546), .Y(ALU_DW01_sub_0__n110) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U141 ( .A(ALU_DW01_sub_0__n548), .Y(ALU_DW01_sub_0__n111) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U142 ( .A(ALU_DW01_sub_0__n652), .Y(ALU_DW01_sub_0__n540) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U143 ( .A(ALU_DW01_sub_0__n403), .Y(ALU_DW01_sub_0__n112) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U144 ( .A(ALU_DW01_sub_0__n391), .Y(ALU_DW01_sub_0__n113) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U145 ( .A(ALU_DW01_sub_0__n393), .Y(ALU_DW01_sub_0__n114) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U146 ( .A(ALU_DW01_sub_0__n400), .Y(ALU_DW01_sub_0__n115) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U147 ( .A(ALU_DW01_sub_0__n404), .Y(ALU_DW01_sub_0__n116) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U148 ( .A(ALU_DW01_sub_0__n394), .Y(ALU_DW01_sub_0__n117) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U149 ( .A(ALU_DW01_sub_0__n396), .Y(ALU_DW01_sub_0__n118) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U150 ( .A(ALU_DW01_sub_0__n474), .Y(ALU_DW01_sub_0__n388) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U151 ( .A(ALU_DW01_sub_0__n376), .Y(ALU_DW01_sub_0__n119) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U152 ( .A(ALU_DW01_sub_0__n699), .Y(ALU_DW01_sub_0__n376) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U153 ( .A(ALU_DW01_sub_0__n713), .Y(ALU_DW01_sub_0__n757) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U154 ( .A(ALU_DW01_sub_0__n288), .Y(ALU_DW01_sub_0__n122) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U155 ( .A(ALU_DW01_sub_0__n408), .Y(ALU_DW01_sub_0__n123) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U156 ( .A(ALU_DW01_sub_0__n420), .Y(ALU_DW01_sub_0__n124) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U157 ( .A(ALU_DW01_sub_0__n126), .Y(ALU_DW01_sub_0__n125) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U158 ( .A(ALU_DW01_sub_0__n769), .Y(ALU_DW01_sub_0__n126) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U159 ( .A(ALU_DW01_sub_0__n306), .Y(ALU__N178) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U160 ( .A(ALU_DW01_sub_0__n136), .Y(ALU_DW01_sub_0__n779) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U161 ( .A(ALU_DW01_sub_0__n779), .Y(ALU_DW01_sub_0__n128) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U162 ( .A(ALU_DW01_sub_0__n717), .Y(ALU_DW01_sub_0__n761) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U163 ( .A(ALU_DW01_sub_0__n41), .Y(ALU__N172) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U164 ( .A(ALU_DW01_sub_0__n131), .Y(ALU_DW01_sub_0__n130) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U165 ( .A(ALU_DW01_sub_0__n211), .Y(ALU_DW01_sub_0__n131) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U166 ( .A(ALU_DW01_sub_0__n538), .Y(ALU_DW01_sub_0__n132) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U167 ( .A(ALU_DW01_sub_0__n550), .Y(ALU_DW01_sub_0__n133) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U168 ( .A(ALU_DW01_sub_0__n244), .Y(ALU__N165) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U169 ( .A(ALU_DW01_sub_0__n245), .Y(ALU_DW01_sub_0__n244) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U170 ( .A(ALU_DW01_sub_0__n768), .Y(ALU_DW01_sub_0__n245) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U171 ( .A(ALU_DW01_sub_0__n264), .Y(ALU__N163) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U172 ( .A(ALU_DW01_sub_0__n265), .Y(ALU_DW01_sub_0__n264) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U173 ( .A(ALU_DW01_sub_0__n770), .Y(ALU_DW01_sub_0__n265) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U174 ( .A(ALU_DW01_sub_0__n330), .Y(ALU_DW01_sub_0__n135) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U175 ( .A(ALU_DW01_sub_0__n681), .Y(ALU_DW01_sub_0__n330) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U176 ( .A(ALU_DW01_sub_0__n57), .B(ALU_DW01_sub_0__n60), .Y(ALU_DW01_sub_0__n136) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U177 ( .A(ALU_DW01_sub_0__n137), .B(ALU_DW01_sub_0__n139), .Y(ALU_DW01_sub_0__n374) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U178 ( .A(ALU_DW01_sub_0__n200), .B(ALU_DW01_sub_0__n362), .Y(ALU_DW01_sub_0__n361) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U179 ( .A(ALU_DW01_sub_0__n58), .Y(ALU_DW01_sub_0__n137) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U180 ( .A(ALU_DW01_sub_0__n370), .Y(ALU_DW01_sub_0__n138) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U181 ( .A(ALU_DW01_sub_0__n359), .B(ALU_DW01_sub_0__n364), .Y(ALU_DW01_sub_0__n363) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U182 ( .A(ALU_DW01_sub_0__n59), .Y(ALU_DW01_sub_0__n139) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U183 ( .A(ALU_DW01_sub_0__n371), .Y(ALU_DW01_sub_0__n140) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U184 ( .A(ALU_DW01_sub_0__n141), .B(ALU_DW01_sub_0__n143), .Y(ALU_DW01_sub_0__n375) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U185 ( .A(ALU_DW01_sub_0__n360), .B(ALU_DW01_sub_0__n366), .Y(ALU_DW01_sub_0__n365) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U186 ( .A(ALU_DW01_sub_0__n61), .Y(ALU_DW01_sub_0__n141) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U187 ( .A(ALU_DW01_sub_0__n372), .Y(ALU_DW01_sub_0__n142) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U188 ( .A(ALU_DW01_sub_0__n360), .B(ALU_DW01_sub_0__n368), .Y(ALU_DW01_sub_0__n367) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U189 ( .A(ALU_DW01_sub_0__n62), .Y(ALU_DW01_sub_0__n143) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U190 ( .A(ALU_DW01_sub_0__n373), .Y(ALU_DW01_sub_0__n144) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U191 ( .A(ALU_DW01_sub_0__n138), .Y(ALU_DW01_sub_0__n362) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U192 ( .A(ALU_DW01_sub_0__n140), .Y(ALU_DW01_sub_0__n364) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U193 ( .A(ALU_DW01_sub_0__n142), .Y(ALU_DW01_sub_0__n366) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U194 ( .A(ALU_DW01_sub_0__n144), .Y(ALU_DW01_sub_0__n368) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U195 ( .A(ALU_DW01_sub_0__n723), .Y(ALU_DW01_sub_0__n765) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U196 ( .A(ALU_DW01_sub_0__n44), .Y(ALU__N168) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U197 ( .A(ALU_DW01_sub_0__n449), .Y(ALU_DW01_sub_0__n146) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U198 ( .A(ALU_DW01_sub_0__n438), .Y(ALU_DW01_sub_0__n147) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U199 ( .A(ALU_DW01_sub_0__n385), .Y(ALU_DW01_sub_0__n148) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U200 ( .A(ALU_DW01_sub_0__n387), .Y(ALU_DW01_sub_0__n149) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U201 ( .A(ALU_DW01_sub_0__n398), .Y(ALU_DW01_sub_0__n150) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U202 ( .A(ALU_DW01_sub_0__n683), .Y(ALU_DW01_sub_0__n151) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U203 ( .A(ALU_DW01_sub_0__n161), .Y(ALU_DW01_sub_0__n683) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U204 ( .A(ALU_DW01_sub_0__n164), .Y(ALU_DW01_sub_0__n152) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U205 ( .A(ALU_DW01_sub_0__n436), .Y(ALU_DW01_sub_0__n153) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U206 ( .A(ALU_DW01_sub_0__n355), .Y(ALU_DW01_sub_0__n154) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U207 ( .A(ALU_DW01_sub_0__n356), .Y(ALU_DW01_sub_0__n155) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U208 ( .A(ALU_DW01_sub_0__n369), .Y(ALU_DW01_sub_0__n156) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U209 ( .A(ALU_DW01_sub_0__n512), .Y(ALU_DW01_sub_0__n157) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U210 ( .A(ALU_DW01_sub_0__n384), .Y(ALU_DW01_sub_0__n158) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U211 ( .A(ALU_DW01_sub_0__n690), .Y(ALU_DW01_sub_0__n384) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U212 ( .A(ALU_DW01_sub_0__n202), .Y(ALU_DW01_sub_0__n159) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U213 ( .A(ALU_DW01_sub_0__n696), .Y(ALU_DW01_sub_0__n202) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U214 ( .A(ALU_DW01_sub_0__n405), .Y(ALU_DW01_sub_0__n160) );
  INVx13_ASAP7_75t_R ALU___ALU_DW01_sub_0___U215 ( .A(ALU_DW01_sub_0__n160), .Y(ALU_DW01_sub_0__n474) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U216 ( .A(ALU_DW01_sub_0__n688), .Y(ALU_DW01_sub_0__n405) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U217 ( .A(ALU__n794), .Y(ALU_DW01_sub_0__n161) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U218 ( .A(ALU_DW01_sub_0__n497), .Y(ALU_DW01_sub_0__n162) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U219 ( .A(ALU_DW01_sub_0__n695), .Y(ALU_DW01_sub_0__n497) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U220 ( .A(ALU_DW01_sub_0__n526), .Y(ALU_DW01_sub_0__n163) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U221 ( .A(ALU_DW01_sub_0__n188), .Y(ALU_DW01_sub_0__n527) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U222 ( .A(ALU_DW01_sub_0__n527), .Y(ALU_DW01_sub_0__n526) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U223 ( .A(ALU_DW01_sub_0__n693), .Y(ALU_DW01_sub_0__n164) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U224 ( .A(ALU_DW01_sub_0__n152), .Y(ALU_DW01_sub_0__n525) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U225 ( .A(ALU_DW01_sub_0__n311), .Y(ALU_DW01_sub_0__n165) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U226 ( .A(ALU_DW01_sub_0__n323), .Y(ALU_DW01_sub_0__n166) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U227 ( .A(n767), .Y(ALU_DW01_sub_0__n677) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U228 ( .A(ALU_DW01_sub_0__n589), .Y(ALU_DW01_sub_0__n168) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U229 ( .A(ALU_DW01_sub_0__n441), .Y(ALU_DW01_sub_0__n590) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U230 ( .A(ALU_DW01_sub_0__n590), .Y(ALU_DW01_sub_0__n589) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U231 ( .A(ALU_DW01_sub_0__n172), .B(ALU_DW01_sub_0__n103), .Y(ALU_DW01_sub_0__n169) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U232 ( .A(ALU_DW01_sub_0__n472), .B(n1010), .Y(ALU_DW01_sub_0__n452) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U233 ( .A(ALU_DW01_sub_0__n101), .Y(ALU_DW01_sub_0__n170) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U234 ( .A(ALU_DW01_sub_0__n647), .B(n1010), .Y(ALU_DW01_sub_0__n453) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U235 ( .A(ALU_DW01_sub_0__n102), .Y(ALU_DW01_sub_0__n171) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U236 ( .A(ALU_DW01_sub_0__n454), .Y(ALU_DW01_sub_0__n172) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U237 ( .A(ALU_DW01_sub_0__n170), .B(ALU_DW01_sub_0__n171), .Y(ALU_DW01_sub_0__n465) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U238 ( .A(ALU_DW01_sub_0__n647), .B(ALU_DW01_sub_0__n472), .Y(ALU_DW01_sub_0__n454) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U239 ( .A(ALU_DW01_sub_0__n28), .Y(ALU_DW01_sub_0__n173) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U240 ( .A(ALU_DW01_sub_0__n685), .Y(ALU_DW01_sub_0__n174) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U241 ( .A(ALU_DW01_sub_0__n157), .Y(ALU_DW01_sub_0__n657) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U242 ( .A(ALU_DW01_sub_0__n122), .Y(ALU_DW01_sub_0__n512) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U243 ( .A(ALU_DW01_sub_0__n174), .Y(ALU_DW01_sub_0__n575) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U244 ( .A(ALU_DW01_sub_0__n106), .B(ALU_DW01_sub_0__n109), .Y(ALU_DW01_sub_0__n175) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U245 ( .A(ALU_DW01_sub_0__n176), .B(ALU_DW01_sub_0__n178), .Y(ALU_DW01_sub_0__n555) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U246 ( .A(ALU_DW01_sub_0__n259), .B(ALU_DW01_sub_0__n543), .Y(ALU_DW01_sub_0__n542) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U247 ( .A(ALU_DW01_sub_0__n107), .Y(ALU_DW01_sub_0__n176) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U248 ( .A(ALU_DW01_sub_0__n551), .Y(ALU_DW01_sub_0__n177) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U249 ( .A(ALU_DW01_sub_0__n540), .B(ALU_DW01_sub_0__n545), .Y(ALU_DW01_sub_0__n544) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U250 ( .A(ALU_DW01_sub_0__n108), .Y(ALU_DW01_sub_0__n178) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U251 ( .A(ALU_DW01_sub_0__n552), .Y(ALU_DW01_sub_0__n179) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U252 ( .A(ALU_DW01_sub_0__n180), .B(ALU_DW01_sub_0__n182), .Y(ALU_DW01_sub_0__n556) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U253 ( .A(ALU_DW01_sub_0__n541), .B(ALU_DW01_sub_0__n547), .Y(ALU_DW01_sub_0__n546) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U254 ( .A(ALU_DW01_sub_0__n110), .Y(ALU_DW01_sub_0__n180) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U255 ( .A(ALU_DW01_sub_0__n553), .Y(ALU_DW01_sub_0__n181) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U256 ( .A(ALU_DW01_sub_0__n541), .B(ALU_DW01_sub_0__n549), .Y(ALU_DW01_sub_0__n548) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U257 ( .A(ALU_DW01_sub_0__n111), .Y(ALU_DW01_sub_0__n182) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U258 ( .A(ALU_DW01_sub_0__n554), .Y(ALU_DW01_sub_0__n183) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U259 ( .A(ALU_DW01_sub_0__n177), .Y(ALU_DW01_sub_0__n543) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U260 ( .A(ALU_DW01_sub_0__n179), .Y(ALU_DW01_sub_0__n545) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U261 ( .A(ALU_DW01_sub_0__n181), .Y(ALU_DW01_sub_0__n547) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U262 ( .A(ALU_DW01_sub_0__n183), .Y(ALU_DW01_sub_0__n549) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U263 ( .A(ALU_DW01_sub_0__n711), .Y(ALU_DW01_sub_0__n756) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U264 ( .A(ALU_DW01_sub_0__n620), .Y(ALU_DW01_sub_0__n185) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U265 ( .A(ALU_DW01_sub_0__n130), .Y(ALU_DW01_sub_0__n572) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U266 ( .A(ALU_DW01_sub_0__n519), .Y(ALU_DW01_sub_0__n186) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U267 ( .A(n1010), .Y(ALU_DW01_sub_0__n457) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U268 ( .A(ALU_DW01_sub_0__n294), .Y(ALU_DW01_sub_0__n187) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U269 ( .A(ALU_DW01_sub_0__n189), .Y(ALU_DW01_sub_0__n188) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U270 ( .A(ALU_DW01_sub_0__n17), .Y(ALU_DW01_sub_0__n189) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U271 ( .A(ALU_DW01_sub_0__n80), .B(ALU_DW01_sub_0__n83), .Y(ALU_DW01_sub_0__n190) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U272 ( .A(ALU_DW01_sub_0__n191), .B(ALU_DW01_sub_0__n193), .Y(ALU_DW01_sub_0__n425) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U273 ( .A(ALU_DW01_sub_0__n347), .B(ALU_DW01_sub_0__n413), .Y(ALU_DW01_sub_0__n412) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U274 ( .A(ALU_DW01_sub_0__n81), .Y(ALU_DW01_sub_0__n191) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U275 ( .A(ALU_DW01_sub_0__n421), .Y(ALU_DW01_sub_0__n192) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U276 ( .A(ALU_DW01_sub_0__n410), .B(ALU_DW01_sub_0__n415), .Y(ALU_DW01_sub_0__n414) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U277 ( .A(ALU_DW01_sub_0__n82), .Y(ALU_DW01_sub_0__n193) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U278 ( .A(ALU_DW01_sub_0__n422), .Y(ALU_DW01_sub_0__n194) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U279 ( .A(ALU_DW01_sub_0__n195), .B(ALU_DW01_sub_0__n197), .Y(ALU_DW01_sub_0__n426) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U280 ( .A(ALU_DW01_sub_0__n411), .B(ALU_DW01_sub_0__n417), .Y(ALU_DW01_sub_0__n416) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U281 ( .A(ALU_DW01_sub_0__n84), .Y(ALU_DW01_sub_0__n195) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U282 ( .A(ALU_DW01_sub_0__n423), .Y(ALU_DW01_sub_0__n196) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U283 ( .A(ALU_DW01_sub_0__n411), .B(ALU_DW01_sub_0__n419), .Y(ALU_DW01_sub_0__n418) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U284 ( .A(ALU_DW01_sub_0__n85), .Y(ALU_DW01_sub_0__n197) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U285 ( .A(ALU_DW01_sub_0__n424), .Y(ALU_DW01_sub_0__n198) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U286 ( .A(ALU_DW01_sub_0__n192), .Y(ALU_DW01_sub_0__n413) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U287 ( .A(ALU_DW01_sub_0__n194), .Y(ALU_DW01_sub_0__n415) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U288 ( .A(ALU_DW01_sub_0__n196), .Y(ALU_DW01_sub_0__n417) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U289 ( .A(ALU_DW01_sub_0__n198), .Y(ALU_DW01_sub_0__n419) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U290 ( .A(n1174), .Y(ALU_DW01_sub_0__n199) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U291 ( .A(n1174), .Y(ALU_DW01_sub_0__n200) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U292 ( .A(ALU_DW01_sub_0__n606), .Y(ALU_DW01_sub_0__n201) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U293 ( .A(ALU__n731), .Y(ALU_DW01_sub_0__n696) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U294 ( .A(ALU_DW01_sub_0__n204), .Y(ALU_DW01_sub_0__n203) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U295 ( .A(ALU_DW01_sub_0__n773), .Y(ALU_DW01_sub_0__n204) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U296 ( .A(ALU_DW01_sub_0__n562), .Y(ALU_DW01_sub_0__n205) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U297 ( .A(ALU_DW01_sub_0__n561), .Y(ALU_DW01_sub_0__n206) );
  CKINVDCx14_ASAP7_75t_R ALU___ALU_DW01_sub_0___U298 ( .A(ALU_DW01_sub_0__n206), .Y(ALU_DW01_sub_0__n654) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U299 ( .A(ALU_DW01_sub_0__n205), .Y(ALU_DW01_sub_0__n561) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U300 ( .A(ALU_DW01_sub_0__n210), .B(ALU_DW01_sub_0__n156), .Y(ALU_DW01_sub_0__n207) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U301 ( .A(ALU_DW01_sub_0__n514), .B(ALU_DW01_sub_0__n200), .Y(ALU_DW01_sub_0__n355) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U302 ( .A(ALU_DW01_sub_0__n154), .Y(ALU_DW01_sub_0__n208) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U303 ( .A(ALU_DW01_sub_0__n670), .B(ALU_DW01_sub_0__n200), .Y(ALU_DW01_sub_0__n356) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U304 ( .A(ALU_DW01_sub_0__n155), .Y(ALU_DW01_sub_0__n209) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U305 ( .A(ALU_DW01_sub_0__n357), .Y(ALU_DW01_sub_0__n210) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U306 ( .A(ALU_DW01_sub_0__n208), .B(ALU_DW01_sub_0__n209), .Y(ALU_DW01_sub_0__n369) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U307 ( .A(ALU_DW01_sub_0__n670), .B(ALU_DW01_sub_0__n514), .Y(ALU_DW01_sub_0__n357) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U308 ( .A(ALU_DW01_sub_0__n216), .B(ALU_DW01_sub_0__n133), .Y(ALU_DW01_sub_0__n211) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U309 ( .A(ALU_DW01_sub_0__n213), .Y(ALU_DW01_sub_0__n212) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U310 ( .A(ALU_DW01_sub_0__n536), .Y(ALU_DW01_sub_0__n213) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U311 ( .A(ALU_DW01_sub_0__n215), .Y(ALU_DW01_sub_0__n214) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U312 ( .A(ALU_DW01_sub_0__n537), .Y(ALU_DW01_sub_0__n215) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U313 ( .A(ALU_DW01_sub_0__n652), .B(ALU_DW01_sub_0__n557), .Y(ALU_DW01_sub_0__n538) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U314 ( .A(ALU_DW01_sub_0__n132), .Y(ALU_DW01_sub_0__n216) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U315 ( .A(ALU_DW01_sub_0__n212), .B(ALU_DW01_sub_0__n214), .Y(ALU_DW01_sub_0__n550) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U316 ( .A(ALU_DW01_sub_0__n557), .B(ALU_DW01_sub_0__n259), .Y(ALU_DW01_sub_0__n536) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U317 ( .A(ALU_DW01_sub_0__n652), .B(ALU_DW01_sub_0__n259), .Y(ALU_DW01_sub_0__n537) );
  CKINVDCx16_ASAP7_75t_R ALU___ALU_DW01_sub_0___U318 ( .A(ALU_DW01_sub_0__n597), .Y(ALU_DW01_sub_0__n652) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U319 ( .A(ALU_DW01_sub_0__n266), .Y(ALU_DW01_sub_0__n306) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U320 ( .A(ALU_DW01_sub_0__n678), .Y(ALU_DW01_sub_0__n217) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U321 ( .A(ALU_DW01_sub_0__n91), .B(ALU_DW01_sub_0__n94), .Y(ALU_DW01_sub_0__n218) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U322 ( .A(ALU_DW01_sub_0__n219), .B(ALU_DW01_sub_0__n221), .Y(ALU_DW01_sub_0__n495) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U323 ( .A(ALU_DW01_sub_0__n345), .B(ALU_DW01_sub_0__n483), .Y(ALU_DW01_sub_0__n482) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U324 ( .A(ALU_DW01_sub_0__n92), .Y(ALU_DW01_sub_0__n219) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U325 ( .A(ALU_DW01_sub_0__n491), .Y(ALU_DW01_sub_0__n220) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U326 ( .A(ALU_DW01_sub_0__n480), .B(ALU_DW01_sub_0__n485), .Y(ALU_DW01_sub_0__n484) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U327 ( .A(ALU_DW01_sub_0__n93), .Y(ALU_DW01_sub_0__n221) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U328 ( .A(ALU_DW01_sub_0__n492), .Y(ALU_DW01_sub_0__n222) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U329 ( .A(ALU_DW01_sub_0__n223), .B(ALU_DW01_sub_0__n225), .Y(ALU_DW01_sub_0__n496) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U330 ( .A(ALU_DW01_sub_0__n481), .B(ALU_DW01_sub_0__n487), .Y(ALU_DW01_sub_0__n486) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U331 ( .A(ALU_DW01_sub_0__n95), .Y(ALU_DW01_sub_0__n223) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U332 ( .A(ALU_DW01_sub_0__n493), .Y(ALU_DW01_sub_0__n224) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U333 ( .A(ALU_DW01_sub_0__n481), .B(ALU_DW01_sub_0__n489), .Y(ALU_DW01_sub_0__n488) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U334 ( .A(ALU_DW01_sub_0__n96), .Y(ALU_DW01_sub_0__n225) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U335 ( .A(ALU_DW01_sub_0__n494), .Y(ALU_DW01_sub_0__n226) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U336 ( .A(ALU_DW01_sub_0__n89), .Y(ALU__N152) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U337 ( .A(ALU_DW01_sub_0__n220), .Y(ALU_DW01_sub_0__n483) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U338 ( .A(ALU_DW01_sub_0__n222), .Y(ALU_DW01_sub_0__n485) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U339 ( .A(ALU_DW01_sub_0__n224), .Y(ALU_DW01_sub_0__n487) );
  NOR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U340 ( .A(ALU_DW01_sub_0__n565), .B(ALU_DW01_sub_0__n480), .Y(ALU_DW01_sub_0__n493) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U341 ( .A(ALU_DW01_sub_0__n226), .Y(ALU_DW01_sub_0__n489) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U342 ( .A(ALU_DW01_sub_0__n66), .B(ALU_DW01_sub_0__n69), .Y(ALU_DW01_sub_0__n227) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U343 ( .A(ALU_DW01_sub_0__n228), .B(ALU_DW01_sub_0__n230), .Y(ALU_DW01_sub_0__n328) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U344 ( .A(ALU_DW01_sub_0__n278), .B(ALU_DW01_sub_0__n316), .Y(ALU_DW01_sub_0__n315) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U345 ( .A(ALU_DW01_sub_0__n67), .Y(ALU_DW01_sub_0__n228) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U346 ( .A(ALU_DW01_sub_0__n324), .Y(ALU_DW01_sub_0__n229) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U347 ( .A(ALU_DW01_sub_0__n313), .B(ALU_DW01_sub_0__n318), .Y(ALU_DW01_sub_0__n317) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U348 ( .A(ALU_DW01_sub_0__n68), .Y(ALU_DW01_sub_0__n230) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U349 ( .A(ALU_DW01_sub_0__n325), .Y(ALU_DW01_sub_0__n231) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U350 ( .A(ALU_DW01_sub_0__n232), .B(ALU_DW01_sub_0__n234), .Y(ALU_DW01_sub_0__n329) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U351 ( .A(ALU_DW01_sub_0__n314), .B(ALU_DW01_sub_0__n320), .Y(ALU_DW01_sub_0__n319) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U352 ( .A(ALU_DW01_sub_0__n70), .Y(ALU_DW01_sub_0__n232) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U353 ( .A(ALU_DW01_sub_0__n326), .Y(ALU_DW01_sub_0__n233) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U354 ( .A(ALU_DW01_sub_0__n314), .B(ALU_DW01_sub_0__n322), .Y(ALU_DW01_sub_0__n321) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U355 ( .A(ALU_DW01_sub_0__n71), .Y(ALU_DW01_sub_0__n234) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U356 ( .A(ALU_DW01_sub_0__n327), .Y(ALU_DW01_sub_0__n235) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U357 ( .A(ALU_DW01_sub_0__n229), .Y(ALU_DW01_sub_0__n316) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U358 ( .A(ALU_DW01_sub_0__n231), .Y(ALU_DW01_sub_0__n318) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U359 ( .A(ALU_DW01_sub_0__n233), .Y(ALU_DW01_sub_0__n320) );
  NOR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U360 ( .A(ALU_DW01_sub_0__n354), .B(ALU_DW01_sub_0__n313), .Y(ALU_DW01_sub_0__n326) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U361 ( .A(ALU_DW01_sub_0__n235), .Y(ALU_DW01_sub_0__n322) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U362 ( .A(ALU_DW01_sub_0__n715), .Y(ALU_DW01_sub_0__n759) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U363 ( .A(ALU__n902), .Y(ALU_DW01_sub_0__n237) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U364 ( .A(ALU_DW01_sub_0__n435), .Y(ALU_DW01_sub_0__n586) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U365 ( .A(ALU_DW01_sub_0__n153), .Y(ALU_DW01_sub_0__n435) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U366 ( .A(ALU_DW01_sub_0__n239), .Y(ALU_DW01_sub_0__n238) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U367 ( .A(ALU_DW01_sub_0__n513), .Y(ALU_DW01_sub_0__n239) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U368 ( .A(ALU_DW01_sub_0__n241), .Y(ALU_DW01_sub_0__n240) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U369 ( .A(ALU_DW01_sub_0__n185), .Y(ALU_DW01_sub_0__n241) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U370 ( .A(ALU_DW01_sub_0__n243), .Y(ALU_DW01_sub_0__n242) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U371 ( .A(ALU_DW01_sub_0__n146), .Y(ALU_DW01_sub_0__n243) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U372 ( .A(ALU_DW01_sub_0__n247), .Y(ALU_DW01_sub_0__n246) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U373 ( .A(ALU_DW01_sub_0__n772), .Y(ALU_DW01_sub_0__n247) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U374 ( .A(ALU_DW01_sub_0__n253), .B(ALU_DW01_sub_0__n166), .Y(ALU_DW01_sub_0__n248) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U375 ( .A(ALU_DW01_sub_0__n250), .Y(ALU_DW01_sub_0__n249) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U376 ( .A(ALU_DW01_sub_0__n309), .Y(ALU_DW01_sub_0__n250) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U377 ( .A(ALU_DW01_sub_0__n252), .Y(ALU_DW01_sub_0__n251) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U378 ( .A(ALU_DW01_sub_0__n310), .Y(ALU_DW01_sub_0__n252) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U379 ( .A(ALU_DW01_sub_0__n659), .B(ALU_DW01_sub_0__n354), .Y(ALU_DW01_sub_0__n311) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U380 ( .A(ALU_DW01_sub_0__n165), .Y(ALU_DW01_sub_0__n253) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U381 ( .A(ALU_DW01_sub_0__n249), .B(ALU_DW01_sub_0__n251), .Y(ALU_DW01_sub_0__n323) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U382 ( .A(ALU_DW01_sub_0__n354), .B(ALU_DW01_sub_0__n278), .Y(ALU_DW01_sub_0__n309) );
  CKINVDCx20_ASAP7_75t_R ALU___ALU_DW01_sub_0___U383 ( .A(ALU_DW01_sub_0__n135), .Y(ALU_DW01_sub_0__n354) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U384 ( .A(ALU_DW01_sub_0__n659), .B(ALU_DW01_sub_0__n278), .Y(ALU_DW01_sub_0__n310) );
  CKINVDCx16_ASAP7_75t_R ALU___ALU_DW01_sub_0___U385 ( .A(ALU_DW01_sub_0__n163), .Y(ALU_DW01_sub_0__n659) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U386 ( .A(ALU_DW01_sub_0__n257), .B(ALU_DW01_sub_0__n150), .Y(ALU_DW01_sub_0__n254) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U387 ( .A(ALU_DW01_sub_0__n474), .B(ALU_DW01_sub_0__n276), .Y(ALU_DW01_sub_0__n385) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U388 ( .A(ALU_DW01_sub_0__n148), .Y(ALU_DW01_sub_0__n255) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U389 ( .A(ALU_DW01_sub_0__n386), .Y(ALU_DW01_sub_0__n256) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U390 ( .A(ALU_DW01_sub_0__n654), .B(ALU_DW01_sub_0__n474), .Y(ALU_DW01_sub_0__n387) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U391 ( .A(ALU_DW01_sub_0__n149), .Y(ALU_DW01_sub_0__n257) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U392 ( .A(ALU_DW01_sub_0__n255), .B(ALU_DW01_sub_0__n256), .Y(ALU_DW01_sub_0__n398) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U393 ( .A(ALU_DW01_sub_0__n654), .B(ALU_DW01_sub_0__n274), .Y(ALU_DW01_sub_0__n386) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U394 ( .A(ALU__n755), .Y(ALU_DW01_sub_0__n258) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U395 ( .A(ALU__n755), .Y(ALU_DW01_sub_0__n259) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U396 ( .A(ALU_DW01_sub_0__n88), .Y(ALU_DW01_sub_0__n650) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U397 ( .A(ALU_DW01_sub_0__n437), .Y(ALU_DW01_sub_0__n602) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U398 ( .A(ALU_DW01_sub_0__n147), .Y(ALU_DW01_sub_0__n437) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U399 ( .A(ALU_DW01_sub_0__n261), .Y(ALU_DW01_sub_0__n260) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U400 ( .A(ALU_DW01_sub_0__n573), .Y(ALU_DW01_sub_0__n261) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U401 ( .A(ALU_DW01_sub_0__n616), .Y(ALU_DW01_sub_0__n262) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U402 ( .A(ALU_DW01_sub_0__n446), .Y(ALU_DW01_sub_0__n263) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U403 ( .A(ALU_DW01_sub_0__n755), .Y(ALU_DW01_sub_0__n266) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U404 ( .A(n892), .Y(ALU_DW01_sub_0__n267) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U405 ( .A(ALU_DW01_sub_0__n704), .Y(ALU_DW01_sub_0__n268) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U406 ( .A(ALU_DW01_sub_0__n242), .Y(ALU_DW01_sub_0__n665) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U407 ( .A(ALU_DW01_sub_0__n268), .Y(ALU_DW01_sub_0__n632) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U408 ( .A(ALU_DW01_sub_0__n700), .Y(ALU_DW01_sub_0__n269) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U409 ( .A(ALU_DW01_sub_0__n7), .Y(ALU_DW01_sub_0__ALU_DW01_sub_0__n772) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U410 ( .A(ALU_DW01_sub_0__n246), .Y(ALU__N161) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U411 ( .A(ALU_DW01_sub_0__n6), .Y(ALU_DW01_sub_0__n781) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U412 ( .A(ALU_DW01_sub_0__n74), .Y(ALU__N151) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U413 ( .A(ALU_DW01_sub_0__n749), .Y(ALU_DW01_sub_0__n780) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U414 ( .A(ALU_DW01_sub_0__n98), .Y(ALU__N153) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U415 ( .A(n1178), .Y(ALU_DW01_sub_0__n273) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U416 ( .A(n1178), .Y(ALU_DW01_sub_0__n274) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U417 ( .A(n1178), .Y(ALU_DW01_sub_0__n275) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U418 ( .A(n1178), .Y(ALU_DW01_sub_0__n276) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U419 ( .A(ALU_DW01_sub_0__n273), .Y(ALU_DW01_sub_0__n390) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U420 ( .A(ALU__n714), .Y(ALU_DW01_sub_0__n277) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U421 ( .A(ALU__n714), .Y(ALU_DW01_sub_0__n278) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U422 ( .A(ALU_DW01_sub_0__n308), .Y(ALU_DW01_sub_0__n279) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U423 ( .A(ALU_DW01_sub_0__n281), .Y(ALU_DW01_sub_0__n280) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U424 ( .A(ALU_DW01_sub_0__n201), .Y(ALU_DW01_sub_0__n281) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U425 ( .A(ALU_DW01_sub_0__n287), .B(ALU_DW01_sub_0__n105), .Y(ALU_DW01_sub_0__n282) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U426 ( .A(ALU_DW01_sub_0__n284), .Y(ALU_DW01_sub_0__n283) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U427 ( .A(ALU_DW01_sub_0__n476), .Y(ALU_DW01_sub_0__n284) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U428 ( .A(ALU_DW01_sub_0__n286), .Y(ALU_DW01_sub_0__n285) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U429 ( .A(ALU_DW01_sub_0__n477), .Y(ALU_DW01_sub_0__n286) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U430 ( .A(ALU_DW01_sub_0__n672), .B(ALU_DW01_sub_0__n565), .Y(ALU_DW01_sub_0__n478) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U431 ( .A(ALU_DW01_sub_0__n104), .Y(ALU_DW01_sub_0__n287) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U432 ( .A(ALU_DW01_sub_0__n283), .B(ALU_DW01_sub_0__n285), .Y(ALU_DW01_sub_0__n490) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U433 ( .A(ALU_DW01_sub_0__n565), .B(ALU_DW01_sub_0__n345), .Y(ALU_DW01_sub_0__n476) );
  CKINVDCx20_ASAP7_75t_R ALU___ALU_DW01_sub_0___U434 ( .A(ALU_DW01_sub_0__n162), .Y(ALU_DW01_sub_0__n565) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U435 ( .A(ALU_DW01_sub_0__n672), .B(ALU_DW01_sub_0__n345), .Y(ALU_DW01_sub_0__n477) );
  CKINVDCx16_ASAP7_75t_R ALU___ALU_DW01_sub_0___U436 ( .A(ALU_DW01_sub_0__n576), .Y(ALU_DW01_sub_0__n672) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U437 ( .A(ALU_DW01_sub_0__n293), .B(ALU_DW01_sub_0__n124), .Y(ALU_DW01_sub_0__n288) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U438 ( .A(ALU_DW01_sub_0__n290), .Y(ALU_DW01_sub_0__n289) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U439 ( .A(ALU_DW01_sub_0__n406), .Y(ALU_DW01_sub_0__n290) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U440 ( .A(ALU_DW01_sub_0__n292), .Y(ALU_DW01_sub_0__n291) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U441 ( .A(ALU_DW01_sub_0__n407), .Y(ALU_DW01_sub_0__n292) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U442 ( .A(ALU_DW01_sub_0__n658), .B(ALU_DW01_sub_0__n427), .Y(ALU_DW01_sub_0__n408) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U443 ( .A(ALU_DW01_sub_0__n123), .Y(ALU_DW01_sub_0__n293) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U444 ( .A(ALU_DW01_sub_0__n289), .B(ALU_DW01_sub_0__n291), .Y(ALU_DW01_sub_0__n420) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U445 ( .A(ALU_DW01_sub_0__n427), .B(ALU_DW01_sub_0__n347), .Y(ALU_DW01_sub_0__n406) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U446 ( .A(ALU_DW01_sub_0__n658), .B(ALU_DW01_sub_0__n347), .Y(ALU_DW01_sub_0__n407) );
  CKINVDCx16_ASAP7_75t_R ALU___ALU_DW01_sub_0___U447 ( .A(ALU_DW01_sub_0__n615), .Y(ALU_DW01_sub_0__n658) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U448 ( .A(ALU_DW01_sub_0__n703), .Y(ALU_DW01_sub_0__n294) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U449 ( .A(ALU_DW01_sub_0__n187), .Y(ALU_DW01_sub_0__n450) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U450 ( .A(ALU_DW01_sub_0__n238), .Y(ALU_DW01_sub_0__n669) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U451 ( .A(n798), .Y(ALU_DW01_sub_0__n700) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U452 ( .A(ALU_DW01_sub_0__n269), .Y(ALU_DW01_sub_0__n628) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U453 ( .A(ALU_DW01_sub_0__n12), .Y(ALU_DW01_sub_0__n295) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U454 ( .A(n794), .Y(ALU_DW01_sub_0__n678) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U455 ( .A(ALU_DW01_sub_0__n217), .Y(ALU_DW01_sub_0__n296) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U456 ( .A(ALU_DW01_sub_0__n619), .Y(ALU_DW01_sub_0__n661) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U457 ( .A(ALU_DW01_sub_0__n240), .Y(ALU_DW01_sub_0__n619) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U458 ( .A(ALU_DW01_sub_0__n112), .B(ALU_DW01_sub_0__n116), .Y(ALU_DW01_sub_0__n297) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U459 ( .A(ALU_DW01_sub_0__n298), .B(ALU_DW01_sub_0__n300), .Y(ALU_DW01_sub_0__n403) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U460 ( .A(ALU_DW01_sub_0__n274), .B(ALU_DW01_sub_0__n392), .Y(ALU_DW01_sub_0__n391) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U461 ( .A(ALU_DW01_sub_0__n113), .Y(ALU_DW01_sub_0__n298) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U462 ( .A(ALU_DW01_sub_0__n399), .Y(ALU_DW01_sub_0__n299) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U463 ( .A(ALU_DW01_sub_0__n389), .B(ALU_DW01_sub_0__n115), .Y(ALU_DW01_sub_0__n393) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U464 ( .A(ALU_DW01_sub_0__n114), .Y(ALU_DW01_sub_0__n300) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U465 ( .A(ALU_DW01_sub_0__n275), .B(ALU_DW01_sub_0__n388), .Y(ALU_DW01_sub_0__n400) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U466 ( .A(ALU_DW01_sub_0__n301), .B(ALU_DW01_sub_0__n303), .Y(ALU_DW01_sub_0__n404) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U467 ( .A(ALU_DW01_sub_0__n390), .B(ALU_DW01_sub_0__n395), .Y(ALU_DW01_sub_0__n394) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U468 ( .A(ALU_DW01_sub_0__n117), .Y(ALU_DW01_sub_0__n301) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U469 ( .A(ALU_DW01_sub_0__n401), .Y(ALU_DW01_sub_0__n302) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U470 ( .A(ALU_DW01_sub_0__n390), .B(ALU_DW01_sub_0__n397), .Y(ALU_DW01_sub_0__n396) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U471 ( .A(ALU_DW01_sub_0__n118), .Y(ALU_DW01_sub_0__n303) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U472 ( .A(ALU_DW01_sub_0__n402), .Y(ALU_DW01_sub_0__n304) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U473 ( .A(ALU_DW01_sub_0__n299), .Y(ALU_DW01_sub_0__n392) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U474 ( .A(ALU_DW01_sub_0__n302), .Y(ALU_DW01_sub_0__n395) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U475 ( .A(ALU_DW01_sub_0__n304), .Y(ALU_DW01_sub_0__n397) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U476 ( .A(ALU_DW01_sub_0__n1), .Y(ALU_DW01_sub_0__n773) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U477 ( .A(ALU_DW01_sub_0__n203), .Y(ALU__N160) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U478 ( .A(ALU_DW01_sub_0__n709), .Y(ALU_DW01_sub_0__n755) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U479 ( .A(n701), .Y(ALU_DW01_sub_0__n685) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U480 ( .A(ALU_DW01_sub_0__n719), .Y(ALU_DW01_sub_0__n762) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U481 ( .A(ALU_DW01_sub_0__n691), .Y(ALU_DW01_sub_0__n308) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U482 ( .A(ALU_DW01_sub_0__n279), .Y(ALU_DW01_sub_0__n378) );
  INVx5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U483 ( .A(ALU_DW01_sub_0__n354), .Y(ALU_DW01_sub_0__n312) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U484 ( .A(ALU_DW01_sub_0__n277), .Y(ALU_DW01_sub_0__n314) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U485 ( .A(ALU_DW01_sub_0__n659), .B(ALU_DW01_sub_0__n354), .Y(ALU_DW01_sub_0__n324) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U486 ( .A(ALU_DW01_sub_0__n277), .B(ALU_DW01_sub_0__n312), .Y(ALU_DW01_sub_0__n325) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U487 ( .A(ALU_DW01_sub_0__n659), .B(ALU_DW01_sub_0__n312), .Y(ALU_DW01_sub_0__n327) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U488 ( .A(n790), .Y(ALU_DW01_sub_0__n681) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U489 ( .A(ALU_DW01_sub_0__n8), .Y(ALU_DW01_sub_0__n331) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U490 ( .A(ALU_DW01_sub_0__n333), .Y(ALU_DW01_sub_0__n332) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U491 ( .A(ALU_DW01_sub_0__n667), .Y(ALU_DW01_sub_0__n333) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U492 ( .A(ALU__n368), .Y(ALU_DW01_sub_0__n702) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U493 ( .A(ALU_DW01_sub_0__n18), .Y(ALU_DW01_sub_0__n334) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U494 ( .A(ALU_DW01_sub_0__n605), .Y(ALU_DW01_sub_0__n662) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U495 ( .A(ALU_DW01_sub_0__n280), .Y(ALU_DW01_sub_0__n605) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U496 ( .A(n352), .Y(ALU_DW01_sub_0__n676) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U497 ( .A(ALU_DW01_sub_0__n47), .B(ALU_DW01_sub_0__n51), .Y(ALU_DW01_sub_0__n335) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U498 ( .A(ALU_DW01_sub_0__n336), .B(ALU_DW01_sub_0__n338), .Y(ALU_DW01_sub_0__n470) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U499 ( .A(n1010), .B(ALU_DW01_sub_0__n459), .Y(ALU_DW01_sub_0__n458) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U500 ( .A(ALU_DW01_sub_0__n48), .Y(ALU_DW01_sub_0__n336) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U501 ( .A(ALU_DW01_sub_0__n466), .Y(ALU_DW01_sub_0__n337) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U502 ( .A(ALU_DW01_sub_0__n456), .B(ALU_DW01_sub_0__n50), .Y(ALU_DW01_sub_0__n460) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U503 ( .A(ALU_DW01_sub_0__n49), .Y(ALU_DW01_sub_0__n338) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U504 ( .A(n1010), .B(ALU_DW01_sub_0__n455), .Y(ALU_DW01_sub_0__n467) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U505 ( .A(ALU_DW01_sub_0__n339), .B(ALU_DW01_sub_0__n341), .Y(ALU_DW01_sub_0__n471) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U506 ( .A(ALU_DW01_sub_0__n457), .B(ALU_DW01_sub_0__n462), .Y(ALU_DW01_sub_0__n461) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U507 ( .A(ALU_DW01_sub_0__n52), .Y(ALU_DW01_sub_0__n339) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U508 ( .A(ALU_DW01_sub_0__n468), .Y(ALU_DW01_sub_0__n340) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U509 ( .A(ALU_DW01_sub_0__n457), .B(ALU_DW01_sub_0__n464), .Y(ALU_DW01_sub_0__n463) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U510 ( .A(ALU_DW01_sub_0__n53), .Y(ALU_DW01_sub_0__n341) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U511 ( .A(ALU_DW01_sub_0__n469), .Y(ALU_DW01_sub_0__n342) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U512 ( .A(ALU_DW01_sub_0__n337), .Y(ALU_DW01_sub_0__n459) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U513 ( .A(ALU_DW01_sub_0__n340), .Y(ALU_DW01_sub_0__n462) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U514 ( .A(ALU_DW01_sub_0__n342), .Y(ALU_DW01_sub_0__n464) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U515 ( .A(ALU_DW01_sub_0__n4), .Y(ALU_DW01_sub_0__n768) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U516 ( .A(ALU__n685), .Y(ALU_DW01_sub_0__n344) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U517 ( .A(ALU__n685), .Y(ALU_DW01_sub_0__n345) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U518 ( .A(ALU__n709), .Y(ALU_DW01_sub_0__n346) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U519 ( .A(ALU__n709), .Y(ALU_DW01_sub_0__n347) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U520 ( .A(ALU_DW01_sub_0__n350), .Y(ALU_DW01_sub_0__n349) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U521 ( .A(ALU_DW01_sub_0__n86), .Y(ALU_DW01_sub_0__n350) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U522 ( .A(ALU_DW01_sub_0__n689), .Y(ALU_DW01_sub_0__n351) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U523 ( .A(ALU_DW01_sub_0__n686), .Y(ALU_DW01_sub_0__n352) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U524 ( .A(ALU_DW01_sub_0__n248), .Y(ALU_DW01_sub_0__n353) );
  INVx5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U525 ( .A(ALU_DW01_sub_0__n514), .Y(ALU_DW01_sub_0__n358) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U526 ( .A(ALU_DW01_sub_0__n670), .Y(ALU_DW01_sub_0__n359) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U527 ( .A(ALU_DW01_sub_0__n199), .Y(ALU_DW01_sub_0__n360) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U528 ( .A(ALU_DW01_sub_0__n670), .B(ALU_DW01_sub_0__n514), .Y(ALU_DW01_sub_0__n370) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U529 ( .A(ALU_DW01_sub_0__n199), .B(ALU_DW01_sub_0__n358), .Y(ALU_DW01_sub_0__n371) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U530 ( .A(ALU_DW01_sub_0__n514), .B(ALU_DW01_sub_0__n359), .Y(ALU_DW01_sub_0__n372) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U531 ( .A(ALU_DW01_sub_0__n670), .B(ALU_DW01_sub_0__n358), .Y(ALU_DW01_sub_0__n373) );
  CKINVDCx16_ASAP7_75t_R ALU___ALU_DW01_sub_0___U532 ( .A(ALU_DW01_sub_0__n119), .Y(ALU_DW01_sub_0__n514) );
  CKINVDCx14_ASAP7_75t_R ALU___ALU_DW01_sub_0___U533 ( .A(ALU_DW01_sub_0__n168), .Y(ALU_DW01_sub_0__n670) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U534 ( .A(ALU__n783), .Y(ALU_DW01_sub_0__n699) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U535 ( .A(ALU_DW01_sub_0__n27), .Y(ALU_DW01_sub_0__n377) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U536 ( .A(n978), .Y(ALU_DW01_sub_0__n691) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U537 ( .A(ALU_DW01_sub_0__n571), .Y(ALU_DW01_sub_0__n651) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U538 ( .A(ALU_DW01_sub_0__n572), .Y(ALU_DW01_sub_0__n571) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U539 ( .A(ALU_DW01_sub_0__n524), .Y(ALU_DW01_sub_0__n379) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U540 ( .A(ALU_DW01_sub_0__n381), .Y(ALU_DW01_sub_0__n380) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U541 ( .A(ALU_DW01_sub_0__n564), .Y(ALU_DW01_sub_0__n381) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U542 ( .A(ALU_DW01_sub_0__n383), .Y(ALU_DW01_sub_0__n382) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U543 ( .A(ALU_DW01_sub_0__n634), .Y(ALU_DW01_sub_0__n383) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U544 ( .A(n851), .Y(ALU_DW01_sub_0__n690) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U545 ( .A(ALU_DW01_sub_0__n654), .Y(ALU_DW01_sub_0__n389) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U546 ( .A(ALU_DW01_sub_0__n654), .B(ALU_DW01_sub_0__n474), .Y(ALU_DW01_sub_0__n399) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U547 ( .A(ALU_DW01_sub_0__n474), .B(ALU_DW01_sub_0__n389), .Y(ALU_DW01_sub_0__n401) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U548 ( .A(ALU_DW01_sub_0__n654), .B(ALU_DW01_sub_0__n388), .Y(ALU_DW01_sub_0__n402) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U549 ( .A(n1056), .Y(ALU_DW01_sub_0__n688) );
  INVx5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U550 ( .A(ALU_DW01_sub_0__n427), .Y(ALU_DW01_sub_0__n409) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U551 ( .A(ALU_DW01_sub_0__n346), .Y(ALU_DW01_sub_0__n411) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U552 ( .A(ALU_DW01_sub_0__n658), .B(ALU_DW01_sub_0__n427), .Y(ALU_DW01_sub_0__n421) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U553 ( .A(ALU_DW01_sub_0__n346), .B(ALU_DW01_sub_0__n409), .Y(ALU_DW01_sub_0__n422) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U554 ( .A(ALU_DW01_sub_0__n427), .B(ALU_DW01_sub_0__n410), .Y(ALU_DW01_sub_0__n423) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U555 ( .A(ALU_DW01_sub_0__n658), .B(ALU_DW01_sub_0__n409), .Y(ALU_DW01_sub_0__n424) );
  CKINVDCx16_ASAP7_75t_R ALU___ALU_DW01_sub_0___U556 ( .A(ALU_DW01_sub_0__n151), .Y(ALU_DW01_sub_0__n427) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U557 ( .A(ALU_DW01_sub_0__n263), .Y(ALU_DW01_sub_0__n615) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U558 ( .A(ALU_DW01_sub_0__n429), .Y(ALU_DW01_sub_0__n428) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U559 ( .A(ALU_DW01_sub_0__n295), .Y(ALU_DW01_sub_0__n429) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U560 ( .A(ALU_DW01_sub_0__n679), .Y(ALU_DW01_sub_0__n430) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U561 ( .A(ALU_DW01_sub_0__n531), .Y(ALU_DW01_sub_0__n612) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U562 ( .A(ALU_DW01_sub_0__n186), .Y(ALU_DW01_sub_0__n577) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U563 ( .A(ALU_DW01_sub_0__n2), .Y(ALU_DW01_sub_0__n770) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U564 ( .A(ALU_DW01_sub_0__n13), .Y(ALU_DW01_sub_0__n432) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U565 ( .A(ALU_DW01_sub_0__n434), .Y(ALU_DW01_sub_0__n433) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U566 ( .A(ALU_DW01_sub_0__n650), .Y(ALU_DW01_sub_0__n434) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U567 ( .A(ALU__n410), .Y(ALU_DW01_sub_0__n692) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U568 ( .A(ALU_DW01_sub_0__n473), .Y(ALU_DW01_sub_0__n653) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U569 ( .A(ALU_DW01_sub_0__n9), .Y(ALU_DW01_sub_0__n436) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U570 ( .A(ALU_DW01_sub_0__n260), .Y(ALU_DW01_sub_0__n656) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U571 ( .A(n1075), .Y(ALU_DW01_sub_0__n686) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U572 ( .A(ALU_DW01_sub_0__n352), .Y(ALU_DW01_sub_0__n588) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U573 ( .A(ALU_DW01_sub_0__n20), .Y(ALU_DW01_sub_0__n438) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U574 ( .A(ALU_DW01_sub_0__n440), .Y(ALU_DW01_sub_0__n439) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U575 ( .A(ALU_DW01_sub_0__n428), .Y(ALU_DW01_sub_0__n440) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U576 ( .A(ALU_DW01_sub_0__n430), .Y(ALU_DW01_sub_0__n604) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U577 ( .A(n1222), .Y(ALU_DW01_sub_0__n679) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U578 ( .A(ALU_DW01_sub_0__n622), .Y(ALU_DW01_sub_0__n663) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U579 ( .A(ALU__n80), .Y(ALU_DW01_sub_0__n675) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U580 ( .A(ALU_DW01_sub_0__n442), .Y(ALU_DW01_sub_0__n441) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U581 ( .A(ALU_DW01_sub_0__n26), .Y(ALU_DW01_sub_0__n442) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U582 ( .A(ALU_DW01_sub_0__n698), .Y(ALU_DW01_sub_0__n443) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U583 ( .A(ALU_DW01_sub_0__n380), .Y(ALU_DW01_sub_0__n671) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U584 ( .A(ALU_DW01_sub_0__n445), .Y(ALU_DW01_sub_0__n444) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U585 ( .A(ALU_DW01_sub_0__n643), .Y(ALU_DW01_sub_0__n445) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U586 ( .A(ALU_DW01_sub_0__n447), .Y(ALU_DW01_sub_0__n446) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U587 ( .A(ALU_DW01_sub_0__n262), .Y(ALU_DW01_sub_0__n447) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U588 ( .A(ALU_DW01_sub_0__n21), .Y(ALU_DW01_sub_0__n449) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U589 ( .A(n619), .Y(ALU_DW01_sub_0__n703) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U590 ( .A(ALU_DW01_sub_0__n633), .Y(ALU_DW01_sub_0__n666) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U591 ( .A(ALU_DW01_sub_0__n382), .Y(ALU_DW01_sub_0__n633) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U592 ( .A(ALU_DW01_sub_0__n725), .Y(ALU_DW01_sub_0__n767) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U593 ( .A(ALU_DW01_sub_0__n54), .Y(ALU__N166) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U594 ( .A(ALU_DW01_sub_0__n647), .Y(ALU_DW01_sub_0__n456) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U595 ( .A(ALU_DW01_sub_0__n647), .B(ALU_DW01_sub_0__n472), .Y(ALU_DW01_sub_0__n466) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U596 ( .A(ALU_DW01_sub_0__n472), .B(ALU_DW01_sub_0__n456), .Y(ALU_DW01_sub_0__n468) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U597 ( .A(ALU_DW01_sub_0__n647), .B(ALU_DW01_sub_0__n455), .Y(ALU_DW01_sub_0__n469) );
  CKINVDCx16_ASAP7_75t_R ALU___ALU_DW01_sub_0___U598 ( .A(ALU_DW01_sub_0__n159), .Y(ALU_DW01_sub_0__n472) );
  CKINVDCx14_ASAP7_75t_R ALU___ALU_DW01_sub_0___U599 ( .A(ALU_DW01_sub_0__n611), .Y(ALU_DW01_sub_0__n647) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U600 ( .A(ALU_DW01_sub_0__n612), .Y(ALU_DW01_sub_0__n611) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U601 ( .A(ALU_DW01_sub_0__n254), .Y(ALU_DW01_sub_0__n473) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U602 ( .A(ALU_DW01_sub_0__n509), .Y(ALU_DW01_sub_0__n475) );
  INVx5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U603 ( .A(ALU_DW01_sub_0__n565), .Y(ALU_DW01_sub_0__n479) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U604 ( .A(ALU_DW01_sub_0__n344), .Y(ALU_DW01_sub_0__n481) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U605 ( .A(ALU_DW01_sub_0__n672), .B(ALU_DW01_sub_0__n565), .Y(ALU_DW01_sub_0__n491) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U606 ( .A(ALU_DW01_sub_0__n344), .B(ALU_DW01_sub_0__n479), .Y(ALU_DW01_sub_0__n492) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U607 ( .A(ALU_DW01_sub_0__n672), .B(ALU_DW01_sub_0__n479), .Y(ALU_DW01_sub_0__n494) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U608 ( .A(ALU_DW01_sub_0__n577), .Y(ALU_DW01_sub_0__n576) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U609 ( .A(ALU__n505), .Y(ALU_DW01_sub_0__n695) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U610 ( .A(ALU_DW01_sub_0__n499), .Y(ALU_DW01_sub_0__n498) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U611 ( .A(ALU_DW01_sub_0__n570), .Y(ALU_DW01_sub_0__n499) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U612 ( .A(ALU_DW01_sub_0__n3), .Y(ALU_DW01_sub_0__n769) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_sub_0___U613 ( .A(ALU_DW01_sub_0__n125), .Y(ALU__N164) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U614 ( .A(ALU_DW01_sub_0__n745), .Y(ALU_DW01_sub_0__n777) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U615 ( .A(ALU_DW01_sub_0__n379), .Y(ALU_DW01_sub_0__n648) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U616 ( .A(ALU_DW01_sub_0__n503), .Y(ALU_DW01_sub_0__n502) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U617 ( .A(ALU_DW01_sub_0__n23), .Y(ALU_DW01_sub_0__n503) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U618 ( .A(ALU_DW01_sub_0__n505), .Y(ALU_DW01_sub_0__n504) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U619 ( .A(ALU_DW01_sub_0__n653), .Y(ALU_DW01_sub_0__n505) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U620 ( .A(ALU_DW01_sub_0__n351), .Y(ALU_DW01_sub_0__n600) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U621 ( .A(n955), .Y(ALU_DW01_sub_0__n689) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U622 ( .A(ALU_DW01_sub_0__n518), .Y(ALU_DW01_sub_0__n506) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U623 ( .A(ALU_DW01_sub_0__n508), .Y(ALU_DW01_sub_0__n507) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U624 ( .A(ALU_DW01_sub_0__n334), .Y(ALU_DW01_sub_0__n508) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U625 ( .A(ALU_DW01_sub_0__n674), .Y(ALU_DW01_sub_0__n509) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U626 ( .A(ALU_DW01_sub_0__n475), .Y(ALU_DW01_sub_0__n624) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U627 ( .A(ALU_DW01_sub_0__n511), .Y(ALU_DW01_sub_0__n510) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U628 ( .A(ALU_DW01_sub_0__n578), .Y(ALU_DW01_sub_0__n511) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U629 ( .A(ALU_DW01_sub_0__n207), .Y(ALU_DW01_sub_0__n513) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U630 ( .A(ALU_DW01_sub_0__n630), .Y(ALU_DW01_sub_0__n515) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U631 ( .A(ALU_DW01_sub_0__n626), .Y(ALU_DW01_sub_0__n516) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U632 ( .A(ALU_DW01_sub_0__n498), .Y(ALU_DW01_sub_0__n646) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U633 ( .A(ALU_DW01_sub_0__n598), .Y(ALU_DW01_sub_0__n517) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U634 ( .A(ALU_DW01_sub_0__n687), .Y(ALU_DW01_sub_0__n518) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U635 ( .A(ALU_DW01_sub_0__n506), .Y(ALU_DW01_sub_0__n563) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U636 ( .A(ALU_DW01_sub_0__n520), .Y(ALU_DW01_sub_0__n519) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U637 ( .A(ALU_DW01_sub_0__n16), .Y(ALU_DW01_sub_0__n520) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U638 ( .A(ALU_DW01_sub_0__n522), .Y(ALU_DW01_sub_0__n521) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U639 ( .A(ALU_DW01_sub_0__n510), .Y(ALU_DW01_sub_0__n522) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U640 ( .A(ALU_DW01_sub_0__n684), .Y(ALU_DW01_sub_0__n523) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U641 ( .A(ALU_DW01_sub_0__n267), .Y(ALU_DW01_sub_0__n673) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U642 ( .A(ALU_DW01_sub_0__n25), .Y(ALU_DW01_sub_0__n524) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U643 ( .A(n1033), .Y(ALU_DW01_sub_0__n693) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U644 ( .A(ALU_DW01_sub_0__n642), .Y(ALU_DW01_sub_0__n649) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U645 ( .A(ALU_DW01_sub_0__n444), .Y(ALU_DW01_sub_0__n642) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U646 ( .A(ALU_DW01_sub_0__n601), .Y(ALU_DW01_sub_0__n660) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U647 ( .A(ALU_DW01_sub_0__n602), .Y(ALU_DW01_sub_0__n601) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U648 ( .A(n547), .Y(ALU_DW01_sub_0__n680) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U649 ( .A(ALU_DW01_sub_0__n623), .Y(ALU_DW01_sub_0__n528) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U650 ( .A(ALU_DW01_sub_0__n739), .Y(ALU_DW01_sub_0__n774) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U651 ( .A(ALU_DW01_sub_0__n721), .Y(ALU_DW01_sub_0__n763) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U652 ( .A(ALU_DW01_sub_0__n532), .Y(ALU_DW01_sub_0__n531) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U653 ( .A(ALU_DW01_sub_0__n29), .Y(ALU_DW01_sub_0__n532) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U654 ( .A(ALU_DW01_sub_0__n534), .Y(ALU_DW01_sub_0__n533) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U655 ( .A(ALU_DW01_sub_0__n648), .Y(ALU_DW01_sub_0__n534) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U656 ( .A(ALU_DW01_sub_0__n694), .Y(ALU_DW01_sub_0__n535) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U657 ( .A(ALU_DW01_sub_0__n535), .Y(ALU_DW01_sub_0__n614) );
  INVx5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U658 ( .A(ALU_DW01_sub_0__n557), .Y(ALU_DW01_sub_0__n539) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U659 ( .A(ALU_DW01_sub_0__n258), .Y(ALU_DW01_sub_0__n541) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U660 ( .A(ALU_DW01_sub_0__n652), .B(ALU_DW01_sub_0__n557), .Y(ALU_DW01_sub_0__n551) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U661 ( .A(ALU_DW01_sub_0__n258), .B(ALU_DW01_sub_0__n539), .Y(ALU_DW01_sub_0__n552) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U662 ( .A(ALU_DW01_sub_0__n557), .B(ALU_DW01_sub_0__n540), .Y(ALU_DW01_sub_0__n553) );
  NOR2x1p5_ASAP7_75t_R ALU___ALU_DW01_sub_0___U663 ( .A(ALU_DW01_sub_0__n652), .B(ALU_DW01_sub_0__n539), .Y(ALU_DW01_sub_0__n554) );
  CKINVDCx16_ASAP7_75t_R ALU___ALU_DW01_sub_0___U664 ( .A(ALU_DW01_sub_0__n158), .Y(ALU_DW01_sub_0__n557) );
  BUFx16f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U665 ( .A(ALU_DW01_sub_0__n517), .Y(ALU_DW01_sub_0__n597) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U666 ( .A(ALU_DW01_sub_0__n559), .Y(ALU_DW01_sub_0__n558) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U667 ( .A(ALU_DW01_sub_0__n507), .Y(ALU_DW01_sub_0__n559) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U668 ( .A(ALU_DW01_sub_0__n701), .Y(ALU_DW01_sub_0__n560) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U669 ( .A(ALU_DW01_sub_0__n22), .Y(ALU_DW01_sub_0__n562) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U670 ( .A(n1162), .Y(ALU_DW01_sub_0__n687) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U671 ( .A(ALU_DW01_sub_0__n585), .Y(ALU_DW01_sub_0__n655) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U672 ( .A(ALU_DW01_sub_0__n586), .Y(ALU_DW01_sub_0__n585) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U673 ( .A(ALU_DW01_sub_0__n282), .Y(ALU_DW01_sub_0__n564) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U674 ( .A(ALU_DW01_sub_0__n567), .Y(ALU_DW01_sub_0__n566) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U675 ( .A(ALU_DW01_sub_0__n515), .Y(ALU_DW01_sub_0__n567) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U676 ( .A(ALU_DW01_sub_0__n569), .Y(ALU_DW01_sub_0__n568) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U677 ( .A(ALU_DW01_sub_0__n516), .Y(ALU_DW01_sub_0__n569) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U678 ( .A(ALU_DW01_sub_0__n169), .Y(ALU_DW01_sub_0__n570) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U679 ( .A(ALU_DW01_sub_0__n173), .Y(ALU_DW01_sub_0__n573) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U680 ( .A(ALU_DW01_sub_0__n657), .Y(ALU_DW01_sub_0__n574) );
  OR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U681 ( .A(ALU_DW01_sub_0__n673), .B(n964), .Y(ALU_DW01_sub_0__n578) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U682 ( .A(n749), .Y(ALU_DW01_sub_0__n684) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U683 ( .A(ALU_DW01_sub_0__n523), .Y(ALU_DW01_sub_0__n579) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U684 ( .A(ALU_DW01_sub_0__n581), .Y(ALU_DW01_sub_0__n580) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U685 ( .A(ALU_DW01_sub_0__n528), .Y(ALU_DW01_sub_0__n581) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U686 ( .A(n888), .Y(ALU_DW01_sub_0__n697) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U687 ( .A(ALU_DW01_sub_0__n747), .Y(ALU_DW01_sub_0__n778) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U688 ( .A(ALU_DW01_sub_0__n584), .Y(ALU_DW01_sub_0__n583) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U689 ( .A(ALU_DW01_sub_0__n353), .Y(ALU_DW01_sub_0__n584) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U690 ( .A(ALU_DW01_sub_0__n656), .Y(ALU_DW01_sub_0__n587) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U691 ( .A(ALU_DW01_sub_0__n671), .Y(ALU_DW01_sub_0__n591) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U692 ( .A(ALU_DW01_sub_0__n237), .Y(ALU_DW01_sub_0__n698) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U693 ( .A(ALU_DW01_sub_0__n443), .Y(ALU_DW01_sub_0__n592) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U694 ( .A(ALU_DW01_sub_0__n741), .Y(ALU_DW01_sub_0__n775) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U695 ( .A(ALU_DW01_sub_0__n595), .Y(ALU_DW01_sub_0__n594) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U696 ( .A(ALU_DW01_sub_0__n583), .Y(ALU_DW01_sub_0__n595) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U697 ( .A(ALU_DW01_sub_0__n682), .Y(ALU_DW01_sub_0__n596) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U698 ( .A(ALU_DW01_sub_0__n596), .Y(ALU_DW01_sub_0__n618) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U699 ( .A(ALU_DW01_sub_0__n502), .Y(ALU_DW01_sub_0__n598) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U700 ( .A(ALU_DW01_sub_0__n504), .Y(ALU_DW01_sub_0__n599) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U701 ( .A(ALU_DW01_sub_0__n439), .Y(ALU_DW01_sub_0__n603) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U702 ( .A(ALU_DW01_sub_0__n15), .Y(ALU_DW01_sub_0__n606) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U703 ( .A(ALU_DW01_sub_0__n675), .Y(ALU_DW01_sub_0__n607) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U704 ( .A(ALU_DW01_sub_0__n580), .Y(ALU_DW01_sub_0__n622) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U705 ( .A(ALU_DW01_sub_0__n24), .Y(ALU_DW01_sub_0__n608) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U706 ( .A(ALU_DW01_sub_0__n560), .Y(ALU_DW01_sub_0__n609) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U707 ( .A(ALU_DW01_sub_0__n625), .Y(ALU_DW01_sub_0__n668) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U708 ( .A(ALU_DW01_sub_0__n568), .Y(ALU_DW01_sub_0__n625) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U709 ( .A(ALU_DW01_sub_0__n743), .Y(ALU_DW01_sub_0__n776) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U710 ( .A(ALU_DW01_sub_0__n533), .Y(ALU_DW01_sub_0__n613) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U711 ( .A(n1123), .Y(ALU_DW01_sub_0__n694) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U712 ( .A(ALU_DW01_sub_0__n30), .Y(ALU_DW01_sub_0__n616) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U713 ( .A(n858), .Y(ALU_DW01_sub_0__n682) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U714 ( .A(ALU_DW01_sub_0__n19), .Y(ALU_DW01_sub_0__n620) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U715 ( .A(ALU_DW01_sub_0__n558), .Y(ALU_DW01_sub_0__n621) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U716 ( .A(ALU_DW01_sub_0__n11), .Y(ALU_DW01_sub_0__n623) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U717 ( .A(n1164), .Y(ALU_DW01_sub_0__n674) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U718 ( .A(ALU_DW01_sub_0__n629), .Y(ALU_DW01_sub_0__n664) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U719 ( .A(ALU_DW01_sub_0__n566), .Y(ALU_DW01_sub_0__n629) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U720 ( .A(ALU_DW01_sub_0__n10), .Y(ALU_DW01_sub_0__n626) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U721 ( .A(ALU_DW01_sub_0__n669), .Y(ALU_DW01_sub_0__n627) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U722 ( .A(ALU_DW01_sub_0__n14), .Y(ALU_DW01_sub_0__n630) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U723 ( .A(ALU_DW01_sub_0__n665), .Y(ALU_DW01_sub_0__n631) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U724 ( .A(n1208), .Y(ALU_DW01_sub_0__n704) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U725 ( .A(ALU_DW01_sub_0__n331), .Y(ALU_DW01_sub_0__n634) );
  BUFx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U726 ( .A(ALU_DW01_sub_0__n608), .Y(ALU_DW01_sub_0__n667) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U727 ( .A(ALU_DW01_sub_0__n702), .Y(ALU_DW01_sub_0__n636) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U728 ( .A(ALU_DW01_sub_0__n646), .Y(ALU_DW01_sub_0__n637) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_sub_0___U729 ( .A(ALU_DW01_sub_0__n733), .Y(ALU_DW01_sub_0__n771) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_sub_0___U730 ( .A(ALU_DW01_sub_0__n640), .Y(ALU_DW01_sub_0__n782) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U731 ( .A(ALU_DW01_sub_0__n782), .Y(ALU__N150) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U732 ( .A(ALU_DW01_sub_0__n641), .Y(ALU_DW01_sub_0__n640) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U733 ( .A(ALU_DW01_sub_0__n752), .Y(ALU_DW01_sub_0__n641) );
  XOR2x2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U734 ( .A(ALU_DW01_sub_0__n673), .B(n964), .Y(ALU_DW01_sub_0__n752) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_sub_0___U735 ( .A(ALU_DW01_sub_0__n432), .Y(ALU_DW01_sub_0__n643) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_sub_0___U736 ( .A(ALU_DW01_sub_0__n433), .Y(ALU_DW01_sub_0__n644) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_sub_0___U737 ( .A(ALU_DW01_sub_0__n692), .Y(ALU_DW01_sub_0__n645) );

 FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_31 ( .A(ALU_DW01_add_1__n301), .B(n888), .CI(n1091), .SN(ALU_DW01_add_1__n383) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_30 ( .A(ALU_DW01_add_1__n360), .B(ALU__n610), .CI(n1010), .CON(ALU_DW01_add_1__n384), .SN(
        n385) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_29 ( .A(n1215), .B(n1123), .CI(ALU_DW01_add_1__n361), .CON(ALU_DW01_add_1__n386), .SN(
        n387) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_28 ( .A(n920), .B(n1033), .CI(ALU_DW01_add_1__n302), .CON(ALU_DW01_add_1__n388), .SN(
        n389) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_26 ( .A(n1100), .B(n978), .CI(ALU_DW01_add_1__n306), .CON(ALU_DW01_add_1__n390), .SN(
        n391) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_25 ( .A(ALU_DW01_add_1__n363), .B(n851), .CI(ALU__n936), .CON(ALU_DW01_add_1__n392), .SN(
        n393) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_24 ( .A(n1064), .B(n955), .CI(ALU_DW01_add_1__n215), .CON(ALU_DW01_add_1__n394), .SN(
        n395) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_23 ( .A(ALU_DW01_add_1__n201), .B(n1056), .CI(n1178), .CON(ALU_DW01_add_1__n396), .SN(
        n397) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_22 ( .A(n1024), .B(n1162), .CI(ALU_DW01_add_1__n366), .CON(ALU_DW01_add_1__n398), .SN(
        n399) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_21 ( .A(n1075), .B(n1225), .CI(ALU_DW01_add_1__n367), .CON(ALU_DW01_add_1__n400), .SN(
        n401) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_20 ( .A(n1068), .B(n701), .CI(ALU_DW01_add_1__n330), .CON(ALU_DW01_add_1__n402), .SN(
        n403) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_19 ( .A(ALU__n1037), .B(ALU__n657), .CI(ALU_DW01_add_1__n368), .CON(ALU_DW01_add_1__n404), .SN(
        n405) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_18 ( .A(n1182), .B(n858), .CI(ALU_DW01_add_1__n194), .CON(ALU_DW01_add_1__n406), .SN(
        n407) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_17 ( .A(n790), .B(ALU__n968), .CI(ALU_DW01_add_1__n370), .CON(ALU_DW01_add_1__n408), .SN(
        n409) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_16 ( .A(n547), .B(n1073), .CI(ALU_DW01_add_1__n335), .CON(ALU_DW01_add_1__n410), .SN(
        n411) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_15 ( .A(n925), .B(n1222), .CI(ALU_DW01_add_1__n371), .CON(ALU_DW01_add_1__n412), .SN(
        n413) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_14 ( .A(n969), .B(n794), .CI(ALU_DW01_add_1__n372), .CON(ALU_DW01_add_1__n414), .SN(
        n415) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_13 ( .A(n767), .B(n1020), .CI(ALU_DW01_add_1__n373), .CON(ALU_DW01_add_1__n416), .SN(
        n417) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_12 ( .A(n352), .B(n1109), .CI(ALU_DW01_add_1__n355), .CON(ALU_DW01_add_1__n418), .SN(
        n419) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_11 ( .A(ALU_DW01_add_1__n375), .B(ALU__n62), .CI(n1152), .CON(ALU_DW01_add_1__n420), .SN(
        n421) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_10 ( .A(n1164), .B(n1229), .CI(ALU_DW01_add_1__n320), .CON(ALU_DW01_add_1__n422), .SN(
        n423) );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_9 ( .A(n1029), .B(n1208), .CI(ALU_DW01_add_1__n377), .CON(ALU_DW01_add_1__n424), .SN(ALU_DW01_add_1__n425)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_8 ( .A(n929), .B(n619), .CI(ALU_DW01_add_1__n378), .CON(ALU_DW01_add_1__n426), .SN(ALU_DW01_add_1__n427)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_7 ( .A(ALU_DW01_add_1__n358), .B(ALU__n111), .CI(n1114), .CON(ALU_DW01_add_1__n428), .SN(ALU_DW01_add_1__n429)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_6 ( .A(n973), .B(ALU__n51), .CI(ALU_DW01_add_1__n332), .CON(ALU_DW01_add_1__n430), .SN(ALU_DW01_add_1__n431)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_5 ( .A(n798), .B(n1233), .CI(ALU_DW01_add_1__n380), .CON(ALU_DW01_add_1__n432), .SN(ALU_DW01_add_1__n433)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_4 ( .A(ALU_DW01_add_1__n263), .B(ALU__n780), .CI(n1174), .CON(ALU_DW01_add_1__n434), .SN(ALU_DW01_add_1__n435)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_3 ( .A(n1060), .B(ALU__n902), .CI(ALU_DW01_add_1__n381), .CON(ALU_DW01_add_1__n436), .SN(ALU_DW01_add_1__n437)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_2 ( .A(ALU_DW01_add_1__n144), .B(ALU__n1033), .CI(ALU__n504), .CON(ALU_DW01_add_1__n438), .SN(ALU_DW01_add_1__n439)
         );
  FAx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U1_1 ( .A(n1015), .B(n749), .CI(ALU_DW01_add_1__n74), .CON(ALU_DW01_add_1__n440), .SN(ALU_DW01_add_1__n441)
         );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U1 ( .A(ALU_DW01_add_1__n391), .Y(ALU_DW01_add_1__n1) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U2 ( .A(ALU_DW01_add_1__n389), .Y(ALU_DW01_add_1__n2) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U3 ( .A(ALU_DW01_add_1__n433), .Y(ALU_DW01_add_1__n3) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U4 ( .A(ALU_DW01_add_1__ALU_DW01_add_1__n411), .Y(ALU_DW01_add_1__n4) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U5 ( .A(ALU_DW01_add_1__n428), .Y(ALU_DW01_add_1__n5) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U6 ( .A(ALU_DW01_add_1__n396), .Y(ALU_DW01_add_1__n6) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_add_1___U7 ( .A(ALU_DW01_add_1__n119), .Y(ALU_DW01_add_1__n358) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_add_1___U8 ( .A(ALU_DW01_add_1__n90), .Y(ALU_DW01_add_1__n201) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U9 ( .A(ALU_DW01_add_1__n438), .Y(ALU_DW01_add_1__n7) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_add_1___U10 ( .A(ALU_DW01_add_1__n63), .Y(ALU_DW01_add_1__n144) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U11 ( .A(ALU_DW01_add_1__n440), .Y(ALU_DW01_add_1__n8) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U12 ( .A(ALU_DW01_add_1__n412), .Y(ALU_DW01_add_1__n9) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U13 ( .A(ALU_DW01_add_1__n414), .Y(ALU_DW01_add_1__n10) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U14 ( .A(ALU_DW01_add_1__n422), .Y(ALU_DW01_add_1__n11) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U15 ( .A(ALU_DW01_add_1__n416), .Y(ALU_DW01_add_1__n12) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U16 ( .A(ALU_DW01_add_1__n426), .Y(ALU_DW01_add_1__n13) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U17 ( .A(ALU_DW01_add_1__n424), .Y(ALU_DW01_add_1__n14) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U18 ( .A(ALU_DW01_add_1__n398), .Y(ALU_DW01_add_1__n15) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U19 ( .A(ALU_DW01_add_1__n432), .Y(ALU_DW01_add_1__n16) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U20 ( .A(ALU_DW01_add_1__n394), .Y(ALU_DW01_add_1__n17) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U21 ( .A(ALU_DW01_add_1__n430), .Y(ALU_DW01_add_1__n18) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U22 ( .A(ALU_DW01_add_1__n388), .Y(ALU_DW01_add_1__n19) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U23 ( .A(ALU_DW01_add_1__n436), .Y(ALU_DW01_add_1__n20) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U24 ( .A(ALU_DW01_add_1__n390), .Y(ALU_DW01_add_1__n21) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U25 ( .A(ALU_DW01_add_1__n402), .Y(ALU_DW01_add_1__n22) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U26 ( .A(ALU_DW01_add_1__n408), .Y(ALU_DW01_add_1__n23) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U27 ( .A(ALU_DW01_add_1__n418), .Y(ALU_DW01_add_1__n24) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U28 ( .A(ALU_DW01_add_1__n386), .Y(ALU_DW01_add_1__n25) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U29 ( .A(ALU_DW01_add_1__n410), .Y(ALU_DW01_add_1__n26) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U30 ( .A(ALU_DW01_add_1__n406), .Y(ALU_DW01_add_1__n27) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U31 ( .A(ALU_DW01_add_1__n404), .Y(ALU_DW01_add_1__n28) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U32 ( .A(ALU_DW01_add_1__n400), .Y(ALU_DW01_add_1__n29) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U33 ( .A(ALU_DW01_add_1__n434), .Y(ALU_DW01_add_1__n30) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U34 ( .A(ALU_DW01_add_1__n420), .Y(ALU_DW01_add_1__n31) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U35 ( .A(ALU_DW01_add_1__n392), .Y(ALU_DW01_add_1__n32) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U36 ( .A(ALU_DW01_add_1__n384), .Y(ALU_DW01_add_1__n33) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_add_1___U37 ( .A(ALU_DW01_add_1__n152), .Y(ALU_DW01_add_1__n263) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_add_1___U38 ( .A(ALU_DW01_add_1__n318), .Y(ALU_DW01_add_1__n375) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_add_1___U39 ( .A(ALU_DW01_add_1__n213), .Y(ALU_DW01_add_1__n363) );
  INVx4_ASAP7_75t_R ALU___ALU_DW01_add_1___U40 ( .A(ALU_DW01_add_1__n205), .Y(ALU_DW01_add_1__n360) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U41 ( .A(ALU__n335), .Y(ALU_DW01_add_1__n34) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U42 ( .A(ALU_DW01_add_1__n334), .Y(ALU_DW01_add_1__n35) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U43 ( .A(ALU_DW01_add_1__n442), .Y(ALU_DW01_add_1__n36) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U44 ( .A(ALU_DW01_add_1__n158), .Y(ALU_DW01_add_1__n157) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U45 ( .A(ALU_DW01_add_1__n38), .Y(ALU_DW01_add_1__n37) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U46 ( .A(ALU_DW01_add_1__n35), .Y(ALU_DW01_add_1__n38) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U47 ( .A(ALU_DW01_add_1__n193), .Y(ALU_DW01_add_1__n39) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U48 ( .A(ALU_DW01_add_1__n143), .Y(ALU_DW01_add_1__n40) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U49 ( .A(ALU_DW01_add_1__n289), .Y(ALU__N145) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U50 ( .A(ALU_DW01_add_1__n43), .Y(ALU_DW01_add_1__n42) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U51 ( .A(ALU_DW01_add_1__n39), .Y(ALU_DW01_add_1__n43) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U52 ( .A(ALU_DW01_add_1__n118), .Y(ALU_DW01_add_1__n44) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U53 ( .A(ALU_DW01_add_1__n105), .Y(ALU_DW01_add_1__n45) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U54 ( .A(ALU_DW01_add_1__n47), .Y(ALU_DW01_add_1__n46) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U55 ( .A(ALU_DW01_add_1__n40), .Y(ALU_DW01_add_1__n47) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U56 ( .A(ALU_DW01_add_1__n23), .Y(ALU_DW01_add_1__n48) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U57 ( .A(ALU_DW01_add_1__n117), .Y(ALU_DW01_add_1__n191) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U58 ( .A(ALU_DW01_add_1__n44), .Y(ALU_DW01_add_1__n117) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U59 ( .A(ALU_DW01_add_1__n64), .Y(ALU_DW01_add_1__n369) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U60 ( .A(ALU_DW01_add_1__n20), .Y(ALU_DW01_add_1__n49) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U61 ( .A(ALU_DW01_add_1__n142), .Y(ALU_DW01_add_1__n381) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U62 ( .A(ALU_DW01_add_1__n46), .Y(ALU_DW01_add_1__n142) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U63 ( .A(ALU_DW01_add_1__n150), .Y(ALU_DW01_add_1__n50) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U64 ( .A(ALU_DW01_add_1__n87), .Y(ALU_DW01_add_1__n51) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U65 ( .A(ALU_DW01_add_1__n53), .Y(ALU_DW01_add_1__n52) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U66 ( .A(ALU_DW01_add_1__n338), .Y(ALU_DW01_add_1__n53) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U67 ( .A(ALU_DW01_add_1__n351), .Y(ALU_DW01_add_1__n255) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U68 ( .A(ALU_DW01_add_1__n255), .Y(ALU_DW01_add_1__n54) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U69 ( .A(ALU_DW01_add_1__n346), .Y(ALU_DW01_add_1__n55) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U70 ( .A(ALU_DW01_add_1__n257), .Y(ALU_DW01_add_1__n56) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U71 ( .A(ALU_DW01_add_1__n347), .Y(ALU_DW01_add_1__n57) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U72 ( .A(ALU_DW01_add_1__n259), .Y(ALU_DW01_add_1__n58) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U73 ( .A(ALU_DW01_add_1__n60), .Y(ALU_DW01_add_1__n59) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U74 ( .A(ALU_DW01_add_1__n94), .Y(ALU_DW01_add_1__n60) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U75 ( .A(n892), .Y(ALU_DW01_add_1__n101) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U76 ( .A(ALU_DW01_add_1__n28), .Y(ALU_DW01_add_1__n61) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U77 ( .A(ALU_DW01_add_1__n192), .Y(ALU_DW01_add_1__n368) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U78 ( .A(ALU_DW01_add_1__n42), .Y(ALU_DW01_add_1__n192) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U79 ( .A(ALU_DW01_add_1__n446), .Y(ALU_DW01_add_1__n62) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U80 ( .A(ALU_DW01_add_1__n104), .Y(ALU_DW01_add_1__n265) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U81 ( .A(ALU_DW01_add_1__n45), .Y(ALU_DW01_add_1__n104) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U82 ( .A(ALU_DW01_add_1__n86), .Y(ALU_DW01_add_1__n156) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U83 ( .A(ALU_DW01_add_1__n51), .Y(ALU_DW01_add_1__n86) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U84 ( .A(ALU_DW01_add_1__n382), .Y(ALU_DW01_add_1__n63) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U85 ( .A(ALU_DW01_add_1__n48), .Y(ALU_DW01_add_1__n64) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U86 ( .A(ALU_DW01_add_1__n333), .Y(ALU_DW01_add_1__n370) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U87 ( .A(ALU_DW01_add_1__n37), .Y(ALU_DW01_add_1__n333) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U88 ( .A(ALU_DW01_add_1__n129), .Y(ALU_DW01_add_1__n65) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U89 ( .A(ALU_DW01_add_1__n348), .Y(ALU_DW01_add_1__n66) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U90 ( .A(ALU_DW01_add_1__n342), .Y(ALU_DW01_add_1__n67) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U91 ( .A(ALU_DW01_add_1__n69), .Y(ALU_DW01_add_1__n68) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U92 ( .A(ALU_DW01_add_1__n444), .Y(ALU_DW01_add_1__n69) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U93 ( .A(ALU_DW01_add_1__n71), .Y(ALU__N148) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U94 ( .A(ALU_DW01_add_1__n233), .Y(ALU_DW01_add_1__n71) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U95 ( .A(ALU_DW01_add_1__n68), .Y(ALU_DW01_add_1__n233) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U96 ( .A(ALU_DW01_add_1__n73), .Y(ALU_DW01_add_1__n72) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U97 ( .A(ALU_DW01_add_1__n369), .Y(ALU_DW01_add_1__n73) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U98 ( .A(ALU_DW01_add_1__n75), .Y(ALU_DW01_add_1__n74) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U99 ( .A(ALU_DW01_add_1__n59), .Y(ALU_DW01_add_1__n75) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U100 ( .A(n964), .B(ALU_DW01_add_1__n101), .Y(ALU_DW01_add_1__n94) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U101 ( .A(ALU_DW01_add_1__n284), .Y(ALU_DW01_add_1__n76) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U102 ( .A(ALU_DW01_add_1__n78), .Y(ALU_DW01_add_1__n77) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U103 ( .A(ALU_DW01_add_1__n62), .Y(ALU_DW01_add_1__n78) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U104 ( .A(ALU_DW01_add_1__n189), .Y(ALU__N146) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U105 ( .A(ALU_DW01_add_1__n81), .Y(ALU_DW01_add_1__n80) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U106 ( .A(ALU_DW01_add_1__n467), .Y(ALU_DW01_add_1__n81) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U107 ( .A(ALU_DW01_add_1__n83), .Y(ALU__N124) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U108 ( .A(ALU_DW01_add_1__n235), .Y(ALU_DW01_add_1__n83) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U109 ( .A(ALU_DW01_add_1__n80), .Y(ALU_DW01_add_1__n235) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U110 ( .A(ALU_DW01_add_1__n85), .Y(ALU_DW01_add_1__n84) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U111 ( .A(ALU_DW01_add_1__n65), .Y(ALU_DW01_add_1__n85) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U112 ( .A(ALU_DW01_add_1__n10), .Y(ALU_DW01_add_1__n87) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U113 ( .A(ALU_DW01_add_1__n33), .Y(ALU_DW01_add_1__n88) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U114 ( .A(ALU_DW01_add_1__n6), .Y(ALU_DW01_add_1__n89) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U115 ( .A(ALU_DW01_add_1__n91), .Y(ALU_DW01_add_1__n90) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U116 ( .A(ALU_DW01_add_1__n365), .Y(ALU_DW01_add_1__n91) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U117 ( .A(ALU_DW01_add_1__n93), .Y(ALU_DW01_add_1__n92) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U118 ( .A(ALU_DW01_add_1__n8), .Y(ALU_DW01_add_1__n93) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U119 ( .A(ALU_DW01_add_1__n322), .Y(ALU_DW01_add_1__n95) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U120 ( .A(ALU_DW01_add_1__n336), .Y(ALU_DW01_add_1__n96) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U121 ( .A(ALU_DW01_add_1__n137), .Y(ALU_DW01_add_1__n97) );
  CKINVDCx8_ASAP7_75t_R ALU___ALU_DW01_add_1___U122 ( .A(ALU_DW01_add_1__n97), .Y(ALU_DW01_add_1__n352) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U123 ( .A(ALU_DW01_add_1__n362), .Y(ALU_DW01_add_1__n137) );
  CKINVDCx5p33_ASAP7_75t_R ALU___ALU_DW01_add_1___U124 ( .A(ALU_DW01_add_1__n352), .Y(ALU_DW01_add_1__n341) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U125 ( .A(ALU_DW01_add_1__n99), .Y(ALU_DW01_add_1__n98) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U126 ( .A(ALU_DW01_add_1__n188), .Y(ALU_DW01_add_1__n99) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U127 ( .A(n892), .Y(ALU_DW01_add_1__n100) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U128 ( .A(ALU_DW01_add_1__n103), .Y(ALU_DW01_add_1__n102) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U129 ( .A(ALU_DW01_add_1__n61), .Y(ALU_DW01_add_1__n103) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U130 ( .A(ALU_DW01_add_1__n13), .Y(ALU_DW01_add_1__n105) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U131 ( .A(ALU_DW01_add_1__n149), .Y(ALU_DW01_add_1__n206) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U132 ( .A(ALU_DW01_add_1__n50), .Y(ALU_DW01_add_1__n149) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U133 ( .A(ALU_DW01_add_1__n107), .Y(ALU_DW01_add_1__n106) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U134 ( .A(ALU_DW01_add_1__n337), .Y(ALU_DW01_add_1__n107) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U135 ( .A(ALU_DW01_add_1__n350), .Y(ALU_DW01_add_1__n184) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U136 ( .A(ALU_DW01_add_1__n184), .Y(ALU_DW01_add_1__n108) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U137 ( .A(ALU_DW01_add_1__n349), .Y(ALU_DW01_add_1__n109) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U138 ( .A(ALU_DW01_add_1__n345), .Y(ALU_DW01_add_1__n110) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U139 ( .A(ALU_DW01_add_1__n187), .Y(ALU_DW01_add_1__n111) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U140 ( .A(ALU_DW01_add_1__n113), .Y(ALU_DW01_add_1__n112) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U141 ( .A(ALU_DW01_add_1__n95), .Y(ALU_DW01_add_1__n113) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U142 ( .A(ALU_DW01_add_1__n115), .Y(ALU_DW01_add_1__n114) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U143 ( .A(ALU_DW01_add_1__n200), .Y(ALU_DW01_add_1__n115) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U144 ( .A(ALU_DW01_add_1__n11), .Y(ALU_DW01_add_1__ALU_DW01_add_1__n116) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U145 ( .A(ALU_DW01_add_1__n84), .Y(ALU_DW01_add_1__n376) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U146 ( .A(ALU_DW01_add_1__n12), .Y(ALU_DW01_add_1__n118) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U147 ( .A(ALU_DW01_add_1__n120), .Y(ALU_DW01_add_1__n119) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U148 ( .A(ALU_DW01_add_1__n379), .Y(ALU_DW01_add_1__n120) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U149 ( .A(ALU_DW01_add_1__n468), .Y(ALU_DW01_add_1__n121) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U150 ( .A(ALU_DW01_add_1__n354), .Y(ALU_DW01_add_1__n122) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U151 ( .A(ALU_DW01_add_1__n326), .Y(ALU_DW01_add_1__n123) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U152 ( .A(ALU_DW01_add_1__n339), .Y(ALU_DW01_add_1__n124) );
  CKINVDCx5p33_ASAP7_75t_R ALU___ALU_DW01_add_1___U153 ( .A(ALU_DW01_add_1__n231), .Y(ALU_DW01_add_1__n274) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U154 ( .A(ALU_DW01_add_1__n232), .Y(ALU_DW01_add_1__n231) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U155 ( .A(ALU_DW01_add_1__n76), .Y(ALU_DW01_add_1__n305) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U156 ( .A(ALU_DW01_add_1__n138), .Y(ALU_DW01_add_1__n125) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U157 ( .A(ALU_DW01_add_1__n127), .Y(ALU_DW01_add_1__n126) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U158 ( .A(ALU_DW01_add_1__n49), .Y(ALU_DW01_add_1__n127) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U159 ( .A(ALU_DW01_add_1__n9), .Y(ALU_DW01_add_1__n128) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U160 ( .A(ALU_DW01_add_1__n155), .Y(ALU_DW01_add_1__n371) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U161 ( .A(ALU_DW01_add_1__n156), .Y(ALU_DW01_add_1__n155) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U162 ( .A(ALU_DW01_add_1__n14), .Y(ALU_DW01_add_1__n129) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U163 ( .A(ALU_DW01_add_1__n264), .Y(ALU_DW01_add_1__n377) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U164 ( .A(ALU_DW01_add_1__n265), .Y(ALU_DW01_add_1__n264) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U165 ( .A(ALU_DW01_add_1__n357), .Y(ALU_DW01_add_1__n130) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U166 ( .A(ALU_DW01_add_1__n307), .Y(ALU_DW01_add_1__n131) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U167 ( .A(ALU_DW01_add_1__n133), .Y(ALU_DW01_add_1__n132) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U168 ( .A(ALU_DW01_add_1__n121), .Y(ALU_DW01_add_1__n133) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U169 ( .A(ALU_DW01_add_1__n204), .Y(ALU__N123) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U170 ( .A(ALU_DW01_add_1__n136), .Y(ALU_DW01_add_1__n135) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U171 ( .A(ALU_DW01_add_1__n123), .Y(ALU_DW01_add_1__n136) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U172 ( .A(ALU_DW01_add_1__n304), .Y(ALU_DW01_add_1__n362) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U173 ( .A(ALU_DW01_add_1__n305), .Y(ALU_DW01_add_1__n304) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U174 ( .A(ALU_DW01_add_1__n299), .Y(ALU_DW01_add_1__n138) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U175 ( .A(ALU_DW01_add_1__n443), .Y(ALU__N149) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U176 ( .A(ALU_DW01_add_1__n125), .Y(ALU_DW01_add_1__n443) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U177 ( .A(ALU_DW01_add_1__n17), .Y(ALU_DW01_add_1__n139) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U178 ( .A(ALU_DW01_add_1__n114), .Y(ALU_DW01_add_1__n364) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U179 ( .A(ALU_DW01_add_1__n141), .Y(ALU_DW01_add_1__n140) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U180 ( .A(ALU_DW01_add_1__n102), .Y(ALU_DW01_add_1__n141) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U181 ( .A(ALU_DW01_add_1__n7), .Y(ALU_DW01_add_1__n143) );
  BUFx4_ASAP7_75t_R ALU___ALU_DW01_add_1___U182 ( .A(ALU_DW01_add_1__n92), .Y(ALU_DW01_add_1__n382) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U183 ( .A(ALU_DW01_add_1__n146), .Y(ALU_DW01_add_1__n145) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U184 ( .A(ALU_DW01_add_1__n131), .Y(ALU_DW01_add_1__n146) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U185 ( .A(ALU_DW01_add_1__n148), .Y(ALU_DW01_add_1__n147) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U186 ( .A(ALU_DW01_add_1__n214), .Y(ALU_DW01_add_1__n148) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U187 ( .A(ALU_DW01_add_1__n34), .Y(ALU_DW01_add_1__ALU_DW01_add_1__n340) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U188 ( .A(ALU_DW01_add_1__n25), .Y(ALU_DW01_add_1__n150) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U189 ( .A(ALU_DW01_add_1__n30), .Y(ALU_DW01_add_1__n151) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U190 ( .A(ALU_DW01_add_1__n153), .Y(ALU_DW01_add_1__n152) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U191 ( .A(ALU_DW01_add_1__n126), .Y(ALU_DW01_add_1__n153) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U192 ( .A(ALU_DW01_add_1__n15), .Y(ALU_DW01_add_1__ALU_DW01_add_1__n154) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U193 ( .A(ALU_DW01_add_1__n321), .Y(ALU_DW01_add_1__n366) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U194 ( .A(ALU_DW01_add_1__n112), .Y(ALU_DW01_add_1__n321) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U195 ( .A(ALU_DW01_add_1__n190), .Y(ALU_DW01_add_1__n372) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U196 ( .A(ALU_DW01_add_1__n191), .Y(ALU_DW01_add_1__n190) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U197 ( .A(ALU_DW01_add_1__n36), .Y(ALU_DW01_add_1__n158) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U198 ( .A(ALU_DW01_add_1__n157), .Y(ALU__N118) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U199 ( .A(ALU_DW01_add_1__n457), .Y(ALU_DW01_add_1__n159) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U200 ( .A(ALU_DW01_add_1__n161), .Y(ALU_DW01_add_1__n160) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U201 ( .A(ALU_DW01_add_1__n458), .Y(ALU_DW01_add_1__n161) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U202 ( .A(ALU_DW01_add_1__n163), .Y(ALU__N133) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U203 ( .A(ALU_DW01_add_1__n313), .Y(ALU_DW01_add_1__n163) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U204 ( .A(ALU_DW01_add_1__n160), .Y(ALU_DW01_add_1__n313) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U205 ( .A(ALU_DW01_add_1__n165), .Y(ALU_DW01_add_1__n164) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U206 ( .A(ALU_DW01_add_1__n464), .Y(ALU_DW01_add_1__n165) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U207 ( .A(ALU_DW01_add_1__n167), .Y(ALU__N127) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U208 ( .A(ALU_DW01_add_1__n295), .Y(ALU_DW01_add_1__n167) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U209 ( .A(ALU_DW01_add_1__n164), .Y(ALU_DW01_add_1__n295) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U210 ( .A(ALU_DW01_add_1__n169), .Y(ALU_DW01_add_1__n168) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U211 ( .A(ALU_DW01_add_1__n122), .Y(ALU_DW01_add_1__n169) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U212 ( .A(ALU_DW01_add_1__n170), .B(ALU_DW01_add_1__n171), .Y(ALU_DW01_add_1__n348) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U213 ( .A(ALU_DW01_add_1__n274), .B(ALU_DW01_add_1__n317), .Y(ALU_DW01_add_1__n342) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U214 ( .A(ALU_DW01_add_1__n67), .Y(ALU_DW01_add_1__n170) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_1___U215 ( .A(ALU_DW01_add_1__n274), .B(ALU_DW01_add_1__n341), .Y(ALU_DW01_add_1__n343) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U216 ( .A(ALU_DW01_add_1__n343), .Y(ALU_DW01_add_1__n171) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U217 ( .A(ALU_DW01_add_1__n98), .Y(ALU_DW01_add_1__n359) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U218 ( .A(ALU_DW01_add_1__n32), .Y(ALU_DW01_add_1__n172) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U219 ( .A(ALU_DW01_add_1__n147), .Y(ALU_DW01_add_1__n213) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U220 ( .A(ALU_DW01_add_1__n174), .Y(ALU_DW01_add_1__n173) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U221 ( .A(ALU_DW01_add_1__n447), .Y(ALU_DW01_add_1__n174) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U222 ( .A(ALU_DW01_add_1__n202), .Y(ALU__N144) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U223 ( .A(ALU_DW01_add_1__n177), .Y(ALU_DW01_add_1__n176) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U224 ( .A(ALU_DW01_add_1__n453), .Y(ALU_DW01_add_1__n177) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U225 ( .A(ALU_DW01_add_1__n179), .Y(ALU_DW01_add_1__n178) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U226 ( .A(ALU_DW01_add_1__n159), .Y(ALU_DW01_add_1__n179) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U227 ( .A(ALU_DW01_add_1__n203), .Y(ALU__N134) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U228 ( .A(ALU_DW01_add_1__n182), .Y(ALU_DW01_add_1__n181) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U229 ( .A(ALU_DW01_add_1__n262), .Y(ALU_DW01_add_1__n182) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U230 ( .A(ALU_DW01_add_1__n108), .Y(ALU_DW01_add_1__n337) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U231 ( .A(ALU_DW01_add_1__n106), .Y(ALU_DW01_add_1__n183) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U232 ( .A(ALU_DW01_add_1__n185), .B(ALU_DW01_add_1__n186), .Y(ALU_DW01_add_1__n350) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_1___U233 ( .A(ALU_DW01_add_1__n341), .B(ALU_DW01_add_1__n109), .Y(ALU_DW01_add_1__n344) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U234 ( .A(ALU_DW01_add_1__n344), .Y(ALU_DW01_add_1__n185) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_1___U235 ( .A(ALU_DW01_add_1__n274), .B(ALU_DW01_add_1__n317), .Y(ALU_DW01_add_1__n349) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U236 ( .A(ALU_DW01_add_1__n274), .B(ALU_DW01_add_1__n111), .Y(ALU_DW01_add_1__n345) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U237 ( .A(ALU_DW01_add_1__n110), .Y(ALU_DW01_add_1__n186) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U238 ( .A(ALU_DW01_add_1__n352), .B(ALU_DW01_add_1__n34), .Y(ALU_DW01_add_1__n187) );
  INVx6_ASAP7_75t_R ALU___ALU_DW01_add_1___U239 ( .A(ALU_DW01_add_1__n340), .Y(ALU_DW01_add_1__n317) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U240 ( .A(ALU_DW01_add_1__n88), .Y(ALU_DW01_add_1__n188) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U241 ( .A(ALU_DW01_add_1__n206), .Y(ALU_DW01_add_1__n205) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U242 ( .A(ALU_DW01_add_1__n2), .Y(ALU_DW01_add_1__n446) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U243 ( .A(ALU_DW01_add_1__n77), .Y(ALU_DW01_add_1__n189) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U244 ( .A(ALU_DW01_add_1__n353), .Y(ALU_DW01_add_1__n373) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U245 ( .A(ALU_DW01_add_1__n168), .Y(ALU_DW01_add_1__n353) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U246 ( .A(ALU_DW01_add_1__n27), .Y(ALU_DW01_add_1__n193) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U247 ( .A(ALU_DW01_add_1__n72), .Y(ALU_DW01_add_1__n194) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U248 ( .A(ALU_DW01_add_1__n329), .Y(ALU_DW01_add_1__n195) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U249 ( .A(ALU_DW01_add_1__n197), .Y(ALU_DW01_add_1__n196) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U250 ( .A(ALU_DW01_add_1__n465), .Y(ALU_DW01_add_1__n197) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U251 ( .A(ALU_DW01_add_1__n199), .Y(ALU_DW01_add_1__n198) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U252 ( .A(ALU_DW01_add_1__n472), .Y(ALU_DW01_add_1__n199) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U253 ( .A(ALU_DW01_add_1__n89), .Y(ALU_DW01_add_1__n200) );
  BUFx4_ASAP7_75t_R ALU___ALU_DW01_add_1___U254 ( .A(ALU_DW01_add_1__n154), .Y(ALU_DW01_add_1__n365) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U255 ( .A(ALU_DW01_add_1__n1), .Y(ALU_DW01_add_1__n447) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U256 ( .A(ALU_DW01_add_1__n173), .Y(ALU_DW01_add_1__n202) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U257 ( .A(ALU_DW01_add_1__n4), .Y(ALU_DW01_add_1__ALU_DW01_add_1__n457) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U258 ( .A(ALU_DW01_add_1__n178), .Y(ALU_DW01_add_1__n203) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U259 ( .A(ALU_DW01_add_1__n3), .Y(ALU_DW01_add_1__n468) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U260 ( .A(ALU_DW01_add_1__n132), .Y(ALU_DW01_add_1__n204) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U261 ( .A(ALU_DW01_add_1__n325), .Y(ALU_DW01_add_1__n361) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U262 ( .A(ALU_DW01_add_1__n135), .Y(ALU_DW01_add_1__n325) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U263 ( .A(ALU_DW01_add_1__n208), .Y(ALU_DW01_add_1__n207) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U264 ( .A(ALU_DW01_add_1__n452), .Y(ALU_DW01_add_1__n208) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U265 ( .A(ALU_DW01_add_1__n210), .Y(ALU_DW01_add_1__n209) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U266 ( .A(ALU_DW01_add_1__n459), .Y(ALU_DW01_add_1__n210) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U267 ( .A(ALU_DW01_add_1__n212), .Y(ALU_DW01_add_1__n211) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U268 ( .A(ALU_DW01_add_1__n130), .Y(ALU_DW01_add_1__n212) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U269 ( .A(ALU_DW01_add_1__n145), .Y(ALU_DW01_add_1__n374) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U270 ( .A(ALU_DW01_add_1__n139), .Y(ALU_DW01_add_1__n214) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U271 ( .A(ALU_DW01_add_1__n364), .Y(ALU_DW01_add_1__n215) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U272 ( .A(ALU_DW01_add_1__n217), .Y(ALU_DW01_add_1__n216) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U273 ( .A(ALU_DW01_add_1__n128), .Y(ALU_DW01_add_1__n217) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U274 ( .A(ALU_DW01_add_1__n16), .Y(ALU_DW01_add_1__n218) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U275 ( .A(ALU_DW01_add_1__n261), .Y(ALU_DW01_add_1__n380) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U276 ( .A(ALU_DW01_add_1__n181), .Y(ALU_DW01_add_1__n261) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U277 ( .A(ALU_DW01_add_1__n220), .Y(ALU_DW01_add_1__n219) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U278 ( .A(ALU_DW01_add_1__n445), .Y(ALU_DW01_add_1__n220) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U279 ( .A(ALU_DW01_add_1__n222), .Y(ALU_DW01_add_1__n221) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U280 ( .A(ALU_DW01_add_1__n463), .Y(ALU_DW01_add_1__n222) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U281 ( .A(ALU_DW01_add_1__n224), .Y(ALU_DW01_add_1__n223) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U282 ( .A(ALU_DW01_add_1__n470), .Y(ALU_DW01_add_1__n224) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U283 ( .A(ALU_DW01_add_1__n226), .Y(ALU_DW01_add_1__n225) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U284 ( .A(ALU_DW01_add_1__n462), .Y(ALU_DW01_add_1__n226) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U285 ( .A(ALU_DW01_add_1__n228), .Y(ALU_DW01_add_1__n227) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U286 ( .A(ALU_DW01_add_1__n466), .Y(ALU_DW01_add_1__n228) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U287 ( .A(ALU_DW01_add_1__n230), .Y(ALU_DW01_add_1__n229) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U288 ( .A(ALU_DW01_add_1__n195), .Y(ALU_DW01_add_1__n230) );
  BUFx12f_ASAP7_75t_R ALU___ALU_DW01_add_1___U289 ( .A(ALU_DW01_add_1__n124), .Y(ALU_DW01_add_1__n232) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U290 ( .A(ALU_DW01_add_1__n385), .Y(ALU_DW01_add_1__n444) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U291 ( .A(ALU_DW01_add_1__n441), .Y(ALU_DW01_add_1__n472) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U292 ( .A(ALU_DW01_add_1__n198), .Y(ALU__N119) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U293 ( .A(ALU_DW01_add_1__n431), .Y(ALU_DW01_add_1__n467) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U294 ( .A(ALU_DW01_add_1__n237), .Y(ALU_DW01_add_1__n236) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U295 ( .A(ALU_DW01_add_1__n172), .Y(ALU_DW01_add_1__n237) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U296 ( .A(ALU_DW01_add_1__n239), .Y(ALU_DW01_add_1__n238) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U297 ( .A(ALU_DW01_add_1__n460), .Y(ALU_DW01_add_1__n239) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U298 ( .A(ALU_DW01_add_1__n241), .Y(ALU_DW01_add_1__n240) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U299 ( .A(ALU_DW01_add_1__n448), .Y(ALU_DW01_add_1__n241) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U300 ( .A(ALU_DW01_add_1__n243), .Y(ALU_DW01_add_1__n242) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U301 ( .A(ALU_DW01_add_1__n450), .Y(ALU_DW01_add_1__n243) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U302 ( .A(ALU_DW01_add_1__n245), .Y(ALU_DW01_add_1__n244) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U303 ( .A(ALU_DW01_add_1__n451), .Y(ALU_DW01_add_1__n245) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U304 ( .A(ALU_DW01_add_1__n247), .Y(ALU_DW01_add_1__n246) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U305 ( .A(ALU_DW01_add_1__n456), .Y(ALU_DW01_add_1__n247) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U306 ( .A(ALU_DW01_add_1__n249), .Y(ALU_DW01_add_1__n248) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U307 ( .A(ALU_DW01_add_1__n461), .Y(ALU_DW01_add_1__n249) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U308 ( .A(ALU_DW01_add_1__n251), .Y(ALU_DW01_add_1__n250) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U309 ( .A(ALU_DW01_add_1__n454), .Y(ALU_DW01_add_1__n251) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U310 ( .A(ALU_DW01_add_1__n253), .Y(ALU_DW01_add_1__n252) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U311 ( .A(ALU_DW01_add_1__n319), .Y(ALU_DW01_add_1__n253) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U312 ( .A(ALU_DW01_add_1__n54), .Y(ALU_DW01_add_1__n338) );
  INVx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U313 ( .A(ALU_DW01_add_1__n52), .Y(ALU_DW01_add_1__n254) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U314 ( .A(ALU_DW01_add_1__n256), .B(ALU_DW01_add_1__n258), .Y(ALU_DW01_add_1__n351) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U315 ( .A(ALU_DW01_add_1__n317), .B(ALU_DW01_add_1__n56), .Y(ALU_DW01_add_1__n346) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U316 ( .A(ALU_DW01_add_1__n55), .Y(ALU_DW01_add_1__n256) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U317 ( .A(ALU_DW01_add_1__n352), .B(n1160), .Y(ALU_DW01_add_1__n257) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U318 ( .A(ALU_DW01_add_1__n341), .B(ALU_DW01_add_1__n58), .Y(ALU_DW01_add_1__n347) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U319 ( .A(ALU_DW01_add_1__n57), .Y(ALU_DW01_add_1__n258) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U320 ( .A(ALU_DW01_add_1__n34), .B(n1160), .Y(ALU_DW01_add_1__n259) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U321 ( .A(ALU_DW01_add_1__n403), .Y(ALU_DW01_add_1__n453) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U322 ( .A(ALU_DW01_add_1__n176), .Y(ALU__N138) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U323 ( .A(ALU_DW01_add_1__n151), .Y(ALU_DW01_add_1__n262) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U324 ( .A(ALU_DW01_add_1__n356), .Y(ALU_DW01_add_1__n378) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U325 ( .A(ALU_DW01_add_1__n211), .Y(ALU_DW01_add_1__n356) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U326 ( .A(ALU_DW01_add_1__n267), .Y(ALU_DW01_add_1__n266) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U327 ( .A(ALU_DW01_add_1__n327), .Y(ALU_DW01_add_1__n267) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U328 ( .A(ALU_DW01_add_1__n269), .Y(ALU_DW01_add_1__n268) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U329 ( .A(ALU_DW01_add_1__n449), .Y(ALU_DW01_add_1__n269) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U330 ( .A(ALU_DW01_add_1__n271), .Y(ALU_DW01_add_1__n270) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U331 ( .A(ALU_DW01_add_1__n455), .Y(ALU_DW01_add_1__n271) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U332 ( .A(ALU_DW01_add_1__n273), .Y(ALU_DW01_add_1__n272) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U333 ( .A(ALU_DW01_add_1__n469), .Y(ALU_DW01_add_1__n273) );
  BUFx10_ASAP7_75t_R ALU___ALU_DW01_add_1___U334 ( .A(n1160), .Y(ALU_DW01_add_1__n339) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U335 ( .A(ALU_DW01_add_1__n387), .Y(ALU_DW01_add_1__n445) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U336 ( .A(ALU_DW01_add_1__n219), .Y(ALU__N147) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U337 ( .A(ALU_DW01_add_1__n397), .Y(ALU_DW01_add_1__n450) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U338 ( .A(ALU_DW01_add_1__n242), .Y(ALU__N141) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U339 ( .A(ALU_DW01_add_1__n401), .Y(ALU_DW01_add_1__n452) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U340 ( .A(ALU_DW01_add_1__n207), .Y(ALU__N139) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U341 ( .A(ALU_DW01_add_1__n423), .Y(ALU_DW01_add_1__n463) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U342 ( .A(ALU_DW01_add_1__n221), .Y(ALU__N128) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U343 ( .A(ALU_DW01_add_1__n419), .Y(ALU_DW01_add_1__n461) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U344 ( .A(ALU_DW01_add_1__n248), .Y(ALU__N130) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U345 ( .A(ALU_DW01_add_1__n429), .Y(ALU_DW01_add_1__n466) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U346 ( .A(ALU_DW01_add_1__n227), .Y(ALU__N125) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U347 ( .A(ALU_DW01_add_1__n421), .Y(ALU_DW01_add_1__n462) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U348 ( .A(ALU_DW01_add_1__n225), .Y(ALU__N129) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U349 ( .A(ALU_DW01_add_1__n283), .Y(ALU_DW01_add_1__n282) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U350 ( .A(ALU_DW01_add_1__n216), .Y(ALU_DW01_add_1__n283) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U351 ( .A(ALU_DW01_add_1__n21), .Y(ALU_DW01_add_1__n284) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U352 ( .A(ALU_DW01_add_1__n286), .Y(ALU_DW01_add_1__n285) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U353 ( .A(ALU_DW01_add_1__n236), .Y(ALU_DW01_add_1__n286) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U354 ( .A(ALU_DW01_add_1__n288), .Y(ALU_DW01_add_1__n287) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U355 ( .A(ALU_DW01_add_1__n218), .Y(ALU_DW01_add_1__n288) );
  AND2x4_ASAP7_75t_R ALU___ALU_DW01_add_1___U356 ( .A(ALU_DW01_add_1__n183), .B(ALU_DW01_add_1__n254), .Y(ALU_DW01_add_1__n289) );
  BUFx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U357 ( .A(ALU_DW01_add_1__n291), .Y(ALU_DW01_add_1__n290) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U358 ( .A(ALU_DW01_add_1__n471), .Y(ALU_DW01_add_1__n291) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U359 ( .A(ALU_DW01_add_1__n399), .Y(ALU_DW01_add_1__n451) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U360 ( .A(ALU_DW01_add_1__n244), .Y(ALU__N140) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U361 ( .A(ALU_DW01_add_1__n407), .Y(ALU_DW01_add_1__n455) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U362 ( .A(ALU_DW01_add_1__n270), .Y(ALU__N136) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U363 ( .A(ALU_DW01_add_1__n409), .Y(ALU_DW01_add_1__n456) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U364 ( .A(ALU_DW01_add_1__n246), .Y(ALU__N135) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U365 ( .A(ALU_DW01_add_1__n425), .Y(ALU_DW01_add_1__n464) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U366 ( .A(ALU_DW01_add_1__n435), .Y(ALU_DW01_add_1__n469) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U367 ( .A(ALU_DW01_add_1__n272), .Y(ALU__N122) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U368 ( .A(ALU_DW01_add_1__n405), .Y(ALU_DW01_add_1__n454) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U369 ( .A(ALU_DW01_add_1__n250), .Y(ALU__N137) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U370 ( .A(ALU_DW01_add_1__n300), .Y(ALU_DW01_add_1__n299) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U371 ( .A(ALU_DW01_add_1__n383), .Y(ALU_DW01_add_1__n300) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U372 ( .A(ALU_DW01_add_1__n359), .Y(ALU_DW01_add_1__n301) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U373 ( .A(ALU_DW01_add_1__n303), .Y(ALU_DW01_add_1__n302) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U374 ( .A(ALU_DW01_add_1__n266), .Y(ALU_DW01_add_1__n303) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U375 ( .A(ALU_DW01_add_1__n285), .Y(ALU_DW01_add_1__n306) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U376 ( .A(ALU_DW01_add_1__n31), .Y(ALU_DW01_add_1__n307) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U377 ( .A(ALU_DW01_add_1__n252), .Y(ALU_DW01_add_1__n318) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U378 ( .A(ALU_DW01_add_1__n309), .Y(ALU_DW01_add_1__n308) );
  BUFx4f_ASAP7_75t_R ALU___ALU_DW01_add_1___U379 ( .A(ALU_DW01_add_1__n287), .Y(ALU_DW01_add_1__n309) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U380 ( .A(ALU_DW01_add_1__n317), .B(ALU_DW01_add_1__n341), .Y(ALU_DW01_add_1__n336) );
  INVx1_ASAP7_75t_R ALU___ALU_DW01_add_1___U381 ( .A(ALU_DW01_add_1__n96), .Y(ALU_DW01_add_1__n310) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U382 ( .A(ALU_DW01_add_1__n393), .Y(ALU_DW01_add_1__n448) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U383 ( .A(ALU_DW01_add_1__n240), .Y(ALU__N143) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U384 ( .A(ALU_DW01_add_1__n395), .Y(ALU_DW01_add_1__n449) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U385 ( .A(ALU_DW01_add_1__n268), .Y(ALU__N142) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U386 ( .A(ALU_DW01_add_1__n413), .Y(ALU_DW01_add_1__n458) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U387 ( .A(ALU_DW01_add_1__n415), .Y(ALU_DW01_add_1__n459) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U388 ( .A(ALU_DW01_add_1__n209), .Y(ALU__N132) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U389 ( .A(ALU_DW01_add_1__n437), .Y(ALU_DW01_add_1__n470) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U390 ( .A(ALU_DW01_add_1__n223), .Y(ALU__N121) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U391 ( .A(ALU_DW01_add_1__n427), .Y(ALU_DW01_add_1__n465) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U392 ( .A(ALU_DW01_add_1__n196), .Y(ALU__N126) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U393 ( .A(ALU_DW01_add_1__n116), .Y(ALU_DW01_add_1__n319) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U394 ( .A(ALU_DW01_add_1__n376), .Y(ALU_DW01_add_1__n320) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U395 ( .A(ALU_DW01_add_1__n29), .Y(ALU_DW01_add_1__n322) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U396 ( .A(ALU_DW01_add_1__n328), .Y(ALU_DW01_add_1__n367) );
  BUFx6f_ASAP7_75t_R ALU___ALU_DW01_add_1___U397 ( .A(ALU_DW01_add_1__n229), .Y(ALU_DW01_add_1__n328) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U398 ( .A(ALU_DW01_add_1__n439), .Y(ALU_DW01_add_1__n471) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U399 ( .A(ALU_DW01_add_1__n290), .Y(ALU__N120) );
  HB1xp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U400 ( .A(ALU_DW01_add_1__n417), .Y(ALU_DW01_add_1__n460) );
  INVxp67_ASAP7_75t_R ALU___ALU_DW01_add_1___U401 ( .A(ALU_DW01_add_1__n238), .Y(ALU__N131) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U402 ( .A(ALU_DW01_add_1__n19), .Y(ALU_DW01_add_1__n326) );
  AND2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U403 ( .A(ALU_DW01_add_1__n310), .B(ALU_DW01_add_1__n66), .Y(ALU_DW01_add_1__n327) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U404 ( .A(ALU_DW01_add_1__n22), .Y(ALU_DW01_add_1__n329) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U405 ( .A(ALU_DW01_add_1__n140), .Y(ALU_DW01_add_1__n330) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U406 ( .A(ALU_DW01_add_1__n18), .Y(ALU_DW01_add_1__n331) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U407 ( .A(ALU_DW01_add_1__n308), .Y(ALU_DW01_add_1__n332) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U408 ( .A(ALU_DW01_add_1__n26), .Y(ALU_DW01_add_1__n334) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U409 ( .A(ALU_DW01_add_1__n282), .Y(ALU_DW01_add_1__n335) );
  XNOR2x2_ASAP7_75t_R ALU___ALU_DW01_add_1___U410 ( .A(ALU_DW01_add_1__n100), .B(n964), .Y(ALU_DW01_add_1__n442) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U411 ( .A(ALU_DW01_add_1__n24), .Y(ALU_DW01_add_1__n354) );
  INVx3_ASAP7_75t_R ALU___ALU_DW01_add_1___U412 ( .A(ALU_DW01_add_1__n374), .Y(ALU_DW01_add_1__n355) );
  BUFx2_ASAP7_75t_R ALU___ALU_DW01_add_1___U413 ( .A(ALU_DW01_add_1__n5), .Y(ALU_DW01_add_1__n357) );
  BUFx4_ASAP7_75t_R ALU___ALU_DW01_add_1___U414 ( .A(ALU_DW01_add_1__n331), .Y(ALU_DW01_add_1__n379) );

  DHLx3_ASAP7_75t_R ALU___output_data_reg_24_ ( .CLK(ALU__n1634), .D(ALU__n1177), .Q(ALU__n1790) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_25_ ( .CLK(ALU__n1634), .D(ALU__n1085), .Q(ALU__n1789) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_26_ ( .CLK(ALU__n1637), .D(ALU__n1230), .Q(ALU__n1788) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_27_ ( .CLK(ALU__n1637), .D(ALU__n810), .Q(ALU__n1787) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_4_ ( .CLK(ALU__n1629), .D(ALU__n1222), .Q(ALU__n1810) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_0_ ( .CLK(ALU__n1633), .D(ALU__n475), .Q(ALU__n1814) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_31_ ( .CLK(ALU__n1639), .D(ALU__n1189), .Q(ALU__n1783) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_5_ ( .CLK(ALU__n1629), .D(ALU__n1267), .Q(ALU__n1809) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_18_ ( .CLK(ALU__n1635), .D(ALU__n995), .Q(ALU__n1796) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_13_ ( .CLK(ALU__n1635), .D(ALU__n1116), .Q(ALU__n1801) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_10_ ( .CLK(ALU__n1632), .D(ALU__n1218), .Q(ALU__n1804) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_3_ ( .CLK(ALU__n1628), .D(ALU__n1141), .Q(ALU__n1811) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_14_ ( .CLK(ALU__n1633), .D(ALU__n1059), .Q(ALU__n1800) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_20_ ( .CLK(ALU__n1636), .D(ALU__n1112), .Q(ALU__n1794) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_11_ ( .CLK(ALU__n1632), .D(ALU__n1137), .Q(ALU__n1803) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_7_ ( .CLK(ALU__n1630), .D(ALU__n1185), .Q(ALU__n1807) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_15_ ( .CLK(ALU__n1633), .D(ALU__n1181), .Q(ALU__n1799) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_21_ ( .CLK(ALU__n1636), .D(ALU__n833), .Q(ALU__n1793) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_29_ ( .CLK(ALU__n1638), .D(ALU__n1026), .Q(ALU__n1785) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_1_ ( .CLK(ALU__n1636), .D(ALU__n1097), .Q(ALU__n1813) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_2_ ( .CLK(ALU__n1628), .D(ALU__n999), .Q(ALU__n1812) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_6_ ( .CLK(ALU__n1630), .D(ALU__n961), .Q(ALU__n1808) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_23_ ( .CLK(ALU__n1635), .D(ALU__n1133), .Q(ALU__n1791) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_17_ ( .CLK(ALU__n1634), .D(ALU__n1089), .Q(ALU__n1797) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_8_ ( .CLK(ALU__n1631), .D(ALU__n930), .Q(ALU__n1806) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_30_ ( .CLK(ALU__n1639), .D(ALU__n991), .Q(ALU__n1784) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_12_ ( .CLK(ALU__n1636), .D(ALU__n1093), .Q(ALU__n1802) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_9_ ( .CLK(ALU__n1631), .D(ALU__n1145), .Q(ALU__n1805) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_19_ ( .CLK(ALU__n1635), .D(ALU__n894), .Q(ALU__n1795) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_16_ ( .CLK(ALU__n1634), .D(ALU__n1263), .Q(ALU__n1798) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_22_ ( .CLK(ALU__n1633), .D(ALU__n1259), .Q(ALU__n1792) );
  DHLx3_ASAP7_75t_R ALU___output_data_reg_28_ ( .CLK(ALU__n1638), .D(ALU__n1226), .Q(ALU__n1786) );
  HB1xp67_ASAP7_75t_R ALU___U3 ( .A(n67), .Y(ALU__n1318) );
  BUFx4_ASAP7_75t_R ALU___U4 ( .A(n8), .Y(ALU__n1080) );
  HB1xp67_ASAP7_75t_R ALU___U5 ( .A(n22), .Y(ALU__n1081) );
  HB1xp67_ASAP7_75t_R ALU___U6 ( .A(n58), .Y(ALU__n1110) );
  HB1xp67_ASAP7_75t_R ALU___U7 ( .A(n23), .Y(ALU__n1166) );
  BUFx12f_ASAP7_75t_R ALU___U8 ( .A(ALU__n4), .Y(ALU__n1) );
  BUFx6f_ASAP7_75t_R ALU___U9 ( .A(ALU__n16), .Y(ALU__n779) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U10 ( .A(ALU__n744), .Y(ALU__n1604) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U11 ( .A(ALU__n777), .Y(ALU__n1598) );
  BUFx12f_ASAP7_75t_R ALU___U12 ( .A(ALU__n5), .Y(ALU__n2) );
  BUFx12f_ASAP7_75t_R ALU___U13 ( .A(ALU__n778), .Y(ALU__n3) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U14 ( .A(ALU__n3), .Y(ALU__n1599) );
  BUFx12f_ASAP7_75t_R ALU___U15 ( .A(ALU__n746), .Y(ALU__n4) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U16 ( .A(ALU__n1), .Y(ALU__ALU__n1602) );
  BUFx12f_ASAP7_75t_R ALU___U17 ( .A(ALU__n1475), .Y(ALU__n5) );
  BUFx4f_ASAP7_75t_R ALU___U18 ( .A(ALU__n1475), .Y(ALU__n7) );
  INVx2_ASAP7_75t_R ALU___U19 ( .A(ALU__n7), .Y(ALU__n21) );
  BUFx12f_ASAP7_75t_R ALU___U20 ( .A(ALU__n764), .Y(ALU__n1475) );
  BUFx16f_ASAP7_75t_R ALU___U21 ( .A(ALU__n468), .Y(ALU__n8) );
  BUFx12f_ASAP7_75t_R ALU___U22 ( .A(ALU__n468), .Y(ALU__n9) );
  INVx13_ASAP7_75t_R ALU___U23 ( .A(ALU__n31), .Y(ALU__n1567) );
  CKINVDCx8_ASAP7_75t_R ALU___U24 ( .A(ALU__n1567), .Y(ALU__n468) );
  INVx4_ASAP7_75t_R ALU___U25 ( .A(ALU__n1485), .Y(ALU__n1055) );
  BUFx2_ASAP7_75t_R ALU___U26 ( .A(ALU__n380), .Y(ALU__n10) );
  INVx2_ASAP7_75t_R ALU___U27 ( .A(ALU__n1258), .Y(ALU__n11) );
  BUFx16f_ASAP7_75t_R ALU___U28 ( .A(ALU__n1576), .Y(ALU__n12) );
  BUFx6f_ASAP7_75t_R ALU___U29 ( .A(ALU__n1576), .Y(ALU__n13) );
  INVx3_ASAP7_75t_R ALU___U30 ( .A(ALU__n1611), .Y(ALU__n1590) );
  INVx3_ASAP7_75t_R ALU___U31 ( .A(ALU__n1611), .Y(ALU__n1589) );
  INVx2_ASAP7_75t_R ALU___U32 ( .A(ALU__n1296), .Y(ALU__n14) );
  BUFx6f_ASAP7_75t_R ALU___U33 ( .A(ALU__n1379), .Y(ALU__n1577) );
  BUFx12f_ASAP7_75t_R ALU___U34 ( .A(ALU__n17), .Y(ALU__n15) );
  BUFx12f_ASAP7_75t_R ALU___U35 ( .A(ALU__n18), .Y(ALU__n16) );
  BUFx12f_ASAP7_75t_R ALU___U36 ( .A(ALU__n677), .Y(ALU__n17) );
  BUFx12f_ASAP7_75t_R ALU___U37 ( .A(ALU__n677), .Y(ALU__n18) );
  BUFx6f_ASAP7_75t_R ALU___U38 ( .A(ALU__n1340), .Y(ALU__n1477) );
  INVx3_ASAP7_75t_R ALU___U39 ( .A(ALU__n1477), .Y(ALU__n19) );
  BUFx12f_ASAP7_75t_R ALU___U40 ( .A(ALU__n1585), .Y(ALU__n20) );
  BUFx12f_ASAP7_75t_R ALU___U41 ( .A(ALU__n20), .Y(ALU__n1571) );
  BUFx12f_ASAP7_75t_R ALU___U42 ( .A(ALU__n1586), .Y(ALU__n1584) );
  BUFx12f_ASAP7_75t_R ALU___U43 ( .A(ALU__n1582), .Y(ALU__n1380) );
  BUFx12f_ASAP7_75t_R ALU___U44 ( .A(ALU__n8), .Y(ALU__n1582) );
  BUFx12f_ASAP7_75t_R ALU___U45 ( .A(ALU__n24), .Y(ALU__n22) );
  BUFx12f_ASAP7_75t_R ALU___U46 ( .A(ALU__n24), .Y(ALU__n23) );
  INVx13_ASAP7_75t_R ALU___U47 ( .A(ALU__n30), .Y(ALU__n1480) );
  BUFx12f_ASAP7_75t_R ALU___U48 ( .A(ALU__n99), .Y(ALU__n24) );
  INVx13_ASAP7_75t_R ALU___U49 ( .A(ALU__n40), .Y(ALU__n1562) );
  BUFx12f_ASAP7_75t_R ALU___U50 ( .A(ALU__n1612), .Y(ALU__n25) );
  BUFx12f_ASAP7_75t_R ALU___U51 ( .A(ALU__n1612), .Y(ALU__n26) );
  INVx3_ASAP7_75t_R ALU___U52 ( .A(ALU__n850), .Y(ALU__n1476) );
  INVx2_ASAP7_75t_R ALU___U53 ( .A(ALU__n1539), .Y(ALU__n27) );
  BUFx12f_ASAP7_75t_R ALU___U54 ( .A(ALU__n1271), .Y(ALU__n1539) );
  BUFx12f_ASAP7_75t_R ALU___U55 ( .A(ALU__n678), .Y(ALU__n28) );
  BUFx12f_ASAP7_75t_R ALU___U56 ( .A(ALU__n678), .Y(ALU__n29) );
  BUFx16f_ASAP7_75t_R ALU___U57 ( .A(ALU__n1492), .Y(ALU__n30) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U58 ( .A(ALU__n1484), .Y(ALU__n850) );
  BUFx16f_ASAP7_75t_R ALU___U59 ( .A(ALU__n46), .Y(ALU__n31) );
  BUFx12f_ASAP7_75t_R ALU___U60 ( .A(ALU__n1570), .Y(ALU__n46) );
  BUFx12f_ASAP7_75t_R ALU___U61 ( .A(ALU__n34), .Y(ALU__n32) );
  BUFx12f_ASAP7_75t_R ALU___U62 ( .A(ALU__n34), .Y(ALU__n33) );
  BUFx12f_ASAP7_75t_R ALU___U63 ( .A(ALU__n70), .Y(ALU__n34) );
  BUFx16f_ASAP7_75t_R ALU___U64 ( .A(ALU__n774), .Y(ALU__n1547) );
  BUFx16f_ASAP7_75t_R ALU___U65 ( .A(ALU__n1573), .Y(ALU__n35) );
  CKINVDCx8_ASAP7_75t_R ALU___U66 ( .A(ALU__n1564), .Y(ALU__n775) );
  CKINVDCx12_ASAP7_75t_R ALU___U67 ( .A(ALU__n35), .Y(ALU__n1564) );
  CKINVDCx9p33_ASAP7_75t_R ALU___U68 ( .A(ALU__n1562), .Y(ALU__n807) );
  BUFx12f_ASAP7_75t_R ALU___U69 ( .A(ALU__n807), .Y(ALU__n1573) );
  BUFx2_ASAP7_75t_R ALU___U70 ( .A(ALU__n697), .Y(ALU__n36) );
  BUFx12f_ASAP7_75t_R ALU___U71 ( .A(ALU__n39), .Y(ALU__n37) );
  BUFx12f_ASAP7_75t_R ALU___U72 ( .A(ALU__n39), .Y(ALU__n38) );
  BUFx12f_ASAP7_75t_R ALU___U73 ( .A(ALU__n75), .Y(ALU__n39) );
  INVx13_ASAP7_75t_R ALU___U74 ( .A(ALU__n45), .Y(ALU__n1534) );
  BUFx16f_ASAP7_75t_R ALU___U75 ( .A(ALU__n1575), .Y(ALU__n40) );
  BUFx12f_ASAP7_75t_R ALU___U76 ( .A(ALU__n1584), .Y(ALU__n1575) );
  BUFx12f_ASAP7_75t_R ALU___U77 ( .A(ALU__n1255), .Y(ALU__n41) );
  BUFx12f_ASAP7_75t_R ALU___U78 ( .A(ALU__n1255), .Y(ALU__n42) );
  BUFx12f_ASAP7_75t_R ALU___U79 ( .A(ALU__n49), .Y(ALU__n43) );
  BUFx12f_ASAP7_75t_R ALU___U80 ( .A(ALU__n49), .Y(ALU__n44) );
  BUFx16f_ASAP7_75t_R ALU___U81 ( .A(ALU__n1542), .Y(ALU__n45) );
  INVx4_ASAP7_75t_R ALU___U82 ( .A(ALU__n1549), .Y(ALU__n1528) );
  BUFx12f_ASAP7_75t_R ALU___U83 ( .A(ALU__n483), .Y(ALU__n1542) );
  BUFx12f_ASAP7_75t_R ALU___U84 ( .A(ALU__n20), .Y(ALU__n1570) );
  BUFx12f_ASAP7_75t_R ALU___U85 ( .A(ALU__n104), .Y(ALU__n47) );
  BUFx12f_ASAP7_75t_R ALU___U86 ( .A(ALU__n104), .Y(ALU__n48) );
  BUFx12f_ASAP7_75t_R ALU___U87 ( .A(ALU__n467), .Y(ALU__n49) );
  BUFx12f_ASAP7_75t_R ALU___U88 ( .A(ALU__n43), .Y(ALU__n50) );
  BUFx12f_ASAP7_75t_R ALU___U89 ( .A(ALU__n1555), .Y(ALU__n1553) );
  INVx6_ASAP7_75t_R ALU___U90 ( .A(ALU__n1583), .Y(ALU__n1556) );
  BUFx12f_ASAP7_75t_R ALU___U91 ( .A(ALU__n72), .Y(ALU__n51) );
  BUFx12f_ASAP7_75t_R ALU___U92 ( .A(ALU__n1370), .Y(ALU__n52) );
  BUFx12f_ASAP7_75t_R ALU___U93 ( .A(ALU__n1370), .Y(ALU__n53) );
  BUFx12f_ASAP7_75t_R ALU___U94 ( .A(ALU__n400), .Y(ALU__n54) );
  BUFx16f_ASAP7_75t_R ALU___U95 ( .A(ALU__n417), .Y(ALU__n55) );
  BUFx12f_ASAP7_75t_R ALU___U96 ( .A(ALU__n808), .Y(ALU__n417) );
  BUFx16f_ASAP7_75t_R ALU___U97 ( .A(ALU__n431), .Y(ALU__n56) );
  BUFx12f_ASAP7_75t_R ALU___U98 ( .A(ALU__n854), .Y(ALU__n431) );
  BUFx12f_ASAP7_75t_R ALU___U99 ( .A(ALU__n1371), .Y(ALU__n57) );
  BUFx12f_ASAP7_75t_R ALU___U100 ( .A(ALU__n1371), .Y(ALU__n58) );
  BUFx12f_ASAP7_75t_R ALU___U101 ( .A(ALU__n61), .Y(ALU__n59) );
  BUFx12f_ASAP7_75t_R ALU___U102 ( .A(ALU__n61), .Y(ALU__n60) );
  BUFx12f_ASAP7_75t_R ALU___U103 ( .A(ALU__n107), .Y(ALU__n61) );
  CKINVDCx10_ASAP7_75t_R ALU___U104 ( .A(ALU__n1540), .Y(ALU__n1537) );
  INVx4_ASAP7_75t_R ALU___U105 ( .A(ALU__n1580), .Y(ALU__n1558) );
  BUFx12f_ASAP7_75t_R ALU___U106 ( .A(ALU__n12), .Y(ALU__n1580) );
  BUFx12f_ASAP7_75t_R ALU___U107 ( .A(ALU__n79), .Y(ALU__n62) );
  BUFx12f_ASAP7_75t_R ALU___U108 ( .A(ALU__n1015), .Y(ALU__n63) );
  BUFx12f_ASAP7_75t_R ALU___U109 ( .A(ALU__n1015), .Y(ALU__n64) );
  BUFx16f_ASAP7_75t_R ALU___U110 ( .A(ALU__n1607), .Y(ALU__n65) );
  BUFx12f_ASAP7_75t_R ALU___U111 ( .A(ALU__n15), .Y(ALU__n1607) );
  BUFx4f_ASAP7_75t_R ALU___U112 ( .A(ALU__n416), .Y(ALU__n66) );
  BUFx4f_ASAP7_75t_R ALU___U113 ( .A(ALU__n430), .Y(ALU__n67) );
  BUFx12f_ASAP7_75t_R ALU___U114 ( .A(ALU__n1130), .Y(ALU__n68) );
  BUFx12f_ASAP7_75t_R ALU___U115 ( .A(ALU__n1130), .Y(ALU__n69) );
  BUFx12f_ASAP7_75t_R ALU___U116 ( .A(ALU__n1614), .Y(ALU__n70) );
  BUFx2_ASAP7_75t_R ALU___U117 ( .A(ALU__n264), .Y(ALU__n71) );
  BUFx12f_ASAP7_75t_R ALU___U118 ( .A(n148), .Y(ALU__n72) );
  BUFx12f_ASAP7_75t_R ALU___U119 ( .A(n148), .Y(ALU__n73) );
  BUFx2_ASAP7_75t_R ALU___U120 ( .A(ALU__n222), .Y(ALU__n74) );
  BUFx12f_ASAP7_75t_R ALU___U121 ( .A(ALU__n776), .Y(ALU__n75) );
  BUFx2_ASAP7_75t_R ALU___U122 ( .A(ALU__n228), .Y(ALU__n76) );
  BUFx16f_ASAP7_75t_R ALU___U129 ( .A(ALU__n1609), .Y(ALU__n77) );
  BUFx6f_ASAP7_75t_R ALU___U130 ( .A(ALU__n1609), .Y(ALU__n78) );
  INVx3_ASAP7_75t_R ALU___U132 ( .A(ALU__n78), .Y(ALU__n1595) );
  BUFx12f_ASAP7_75t_R ALU___U133 ( .A(n389), .Y(ALU__n79) );
  BUFx12f_ASAP7_75t_R ALU___U136 ( .A(n389), .Y(ALU__n80) );
  BUFx2_ASAP7_75t_R ALU___U137 ( .A(ALU__n168), .Y(ALU__n81) );
  AO22x2_ASAP7_75t_R ALU___U138 ( .A1(ALU__N176), .A2(ALU__n1566), .B1(ALU__N285), .B2(ALU__n1528), .Y(
        n168) );
  BUFx2_ASAP7_75t_R ALU___U139 ( .A(ALU__n192), .Y(ALU__n82) );
  BUFx3_ASAP7_75t_R ALU___U143 ( .A(ALU__n84), .Y(ALU__n83) );
  BUFx2_ASAP7_75t_R ALU___U144 ( .A(ALU__n210), .Y(ALU__n84) );
  AO22x2_ASAP7_75t_R ALU___U145 ( .A1(ALU__N169), .A2(ALU__n1563), .B1(ALU__N278), .B2(ALU__n1533), .Y(
        n210) );
  BUFx4f_ASAP7_75t_R ALU___U146 ( .A(ALU__n83), .Y(ALU__n374) );
  BUFx3_ASAP7_75t_R ALU___U150 ( .A(ALU__n86), .Y(ALU__n85) );
  INVx2_ASAP7_75t_R ALU___U151 ( .A(ALU__n96), .Y(ALU__n86) );
  CKINVDCx14_ASAP7_75t_R ALU___U152 ( .A(ALU__n464), .Y(ALU__n1624) );
  INVx3_ASAP7_75t_R ALU___U153 ( .A(ALU__n612), .Y(ALU__n1469) );
  BUFx3_ASAP7_75t_R ALU___U157 ( .A(ALU__n88), .Y(ALU__n87) );
  BUFx2_ASAP7_75t_R ALU___U158 ( .A(ALU__n162), .Y(ALU__n88) );
  AO22x2_ASAP7_75t_R ALU___U159 ( .A1(ALU__N177), .A2(ALU__n1566), .B1(ALU__N286), .B2(ALU__n1537), .Y(
        n162) );
  BUFx4f_ASAP7_75t_R ALU___U160 ( .A(ALU__n87), .Y(ALU__n95) );
  BUFx2_ASAP7_75t_R ALU___U164 ( .A(ALU__n174), .Y(ALU__n89) );
  BUFx2_ASAP7_75t_R ALU___U165 ( .A(ALU__n216), .Y(ALU__n90) );
  BUFx16f_ASAP7_75t_R ALU___U167 ( .A(ALU__n1625), .Y(ALU__n91) );
  BUFx12f_ASAP7_75t_R ALU___U171 ( .A(ALU__n1295), .Y(ALU__n1625) );
  BUFx12f_ASAP7_75t_R ALU___U172 ( .A(ALU__n115), .Y(ALU__n92) );
  BUFx12f_ASAP7_75t_R ALU___U174 ( .A(ALU__n115), .Y(ALU__n93) );
  BUFx4f_ASAP7_75t_R ALU___U178 ( .A(ALU__n95), .Y(ALU__n94) );
  INVx2_ASAP7_75t_R ALU___U179 ( .A(ALU__n94), .Y(ALU__n837) );
  BUFx12f_ASAP7_75t_R ALU___U181 ( .A(ALU__n103), .Y(ALU__n96) );
  BUFx12f_ASAP7_75t_R ALU___U185 ( .A(ALU__n103), .Y(ALU__n97) );
  BUFx16f_ASAP7_75t_R ALU___U186 ( .A(ALU__n1076), .Y(ALU__n98) );
  CKINVDCx9p33_ASAP7_75t_R ALU___U187 ( .A(ALU__n98), .Y(ALU__n1470) );
  BUFx12f_ASAP7_75t_R ALU___U188 ( .A(ALU__n1078), .Y(ALU__n1076) );
  BUFx12f_ASAP7_75t_R ALU___U192 ( .A(ALU__n1606), .Y(ALU__n99) );
  INVx6_ASAP7_75t_R ALU___U193 ( .A(ALU__n432), .Y(ALU__n1362) );
  BUFx2_ASAP7_75t_R ALU___U195 ( .A(ALU__n180), .Y(ALU__n100) );
  AO22x2_ASAP7_75t_R ALU___U199 ( .A1(ALU__N174), .A2(ALU__n1565), .B1(ALU__N283), .B2(ALU__n1536), .Y(
        n180) );
  BUFx4f_ASAP7_75t_R ALU___U200 ( .A(ALU__n102), .Y(ALU__n101) );
  BUFx3_ASAP7_75t_R ALU___U201 ( .A(ALU__n81), .Y(ALU__n102) );
  BUFx12f_ASAP7_75t_R ALU___U202 ( .A(ALU__n652), .Y(ALU__n103) );
  BUFx12f_ASAP7_75t_R ALU___U206 ( .A(ALU__n1499), .Y(ALU__n104) );
  BUFx12f_ASAP7_75t_R ALU___U207 ( .A(ALU__n60), .Y(ALU__n105) );
  BUFx12f_ASAP7_75t_R ALU___U209 ( .A(ALU__n59), .Y(ALU__n106) );
  BUFx12f_ASAP7_75t_R ALU___U213 ( .A(ALU__n499), .Y(ALU__n107) );
  BUFx2_ASAP7_75t_R ALU___U214 ( .A(ALU__n186), .Y(ALU__n108) );
  BUFx4f_ASAP7_75t_R ALU___U215 ( .A(ALU__n110), .Y(ALU__n109) );
  BUFx3_ASAP7_75t_R ALU___U216 ( .A(ALU__n100), .Y(ALU__n110) );
  BUFx12f_ASAP7_75t_R ALU___U220 ( .A(ALU__n367), .Y(ALU__n111) );
  BUFx16f_ASAP7_75t_R ALU___U221 ( .A(ALU__n650), .Y(ALU__n112) );
  BUFx12f_ASAP7_75t_R ALU___U222 ( .A(ALU__n96), .Y(ALU__n650) );
  BUFx12f_ASAP7_75t_R ALU___U223 ( .A(ALU__n93), .Y(ALU__n113) );
  BUFx12f_ASAP7_75t_R ALU___U227 ( .A(ALU__n92), .Y(ALU__n114) );
  BUFx12f_ASAP7_75t_R ALU___U228 ( .A(ALU__n1491), .Y(ALU__n115) );
  CKINVDCx12_ASAP7_75t_R ALU___U229 ( .A(ALU__n1523), .Y(ALU__n1515) );
  BUFx16f_ASAP7_75t_R ALU___U230 ( .A(ALU__n343), .Y(ALU__n116) );
  BUFx12f_ASAP7_75t_R ALU___U234 ( .A(ALU__n704), .Y(ALU__n343) );
  INVx4_ASAP7_75t_R ALU___U235 ( .A(ALU__n334), .Y(ALU__n1685) );
  BUFx3_ASAP7_75t_R ALU___U236 ( .A(ALU__n134), .Y(ALU__n130) );
  BUFx2_ASAP7_75t_R ALU___U237 ( .A(ALU__n198), .Y(ALU__n134) );
  AO22x2_ASAP7_75t_R ALU___U241 ( .A1(ALU__N171), .A2(ALU__n1563), .B1(ALU__N280), .B2(ALU__n1537), .Y(
        n198) );
  BUFx4f_ASAP7_75t_R ALU___U242 ( .A(ALU__n130), .Y(ALU__n360) );
  BUFx4f_ASAP7_75t_R ALU___U243 ( .A(ALU__n331), .Y(ALU__n138) );
  BUFx3_ASAP7_75t_R ALU___U244 ( .A(ALU__n108), .Y(ALU__n331) );
  BUFx12f_ASAP7_75t_R ALU___U248 ( .A(ALU__n349), .Y(ALU__n332) );
  BUFx12f_ASAP7_75t_R ALU___U249 ( .A(ALU__n349), .Y(ALU__n333) );
  BUFx16f_ASAP7_75t_R ALU___U251 ( .A(ALU__n409), .Y(ALU__n334) );
  BUFx12f_ASAP7_75t_R ALU___U255 ( .A(ALU__n336), .Y(ALU__n335) );
  BUFx12f_ASAP7_75t_R ALU___U256 ( .A(n435), .Y(ALU__n336) );
  BUFx16f_ASAP7_75t_R ALU___U258 ( .A(ALU__n651), .Y(ALU__n337) );
  CKINVDCx9p33_ASAP7_75t_R ALU___U262 ( .A(ALU__n337), .Y(ALU__n1618) );
  BUFx12f_ASAP7_75t_R ALU___U263 ( .A(ALU__n97), .Y(ALU__n651) );
  BUFx4f_ASAP7_75t_R ALU___U265 ( .A(ALU__n339), .Y(ALU__n338) );
  BUFx3_ASAP7_75t_R ALU___U269 ( .A(ALU__n36), .Y(ALU__n339) );
  BUFx2_ASAP7_75t_R ALU___U270 ( .A(ALU__n1398), .Y(ALU__n340) );
  BUFx2_ASAP7_75t_R ALU___U271 ( .A(ALU__n1399), .Y(ALU__n341) );
  OR2x2_ASAP7_75t_R ALU___U272 ( .A(ALU__n1397), .B(ALU__n341), .Y(ALU__n697) );
  OR2x2_ASAP7_75t_R ALU___U276 ( .A(ALU_ctl[0]), .B(ALU__n1406), .Y(ALU__n1399) );
  BUFx2_ASAP7_75t_R ALU___U277 ( .A(ALU__n258), .Y(ALU__n342) );
  BUFx12f_ASAP7_75t_R ALU___U279 ( .A(ALU__n25), .Y(ALU__n704) );
  BUFx4f_ASAP7_75t_R ALU___U283 ( .A(ALU__n345), .Y(ALU__n344) );
  BUFx3_ASAP7_75t_R ALU___U284 ( .A(ALU__n89), .Y(ALU__n345) );
  BUFx4f_ASAP7_75t_R ALU___U286 ( .A(ALU__n347), .Y(ALU__n346) );
  BUFx3_ASAP7_75t_R ALU___U290 ( .A(ALU__n82), .Y(ALU__n347) );
  AO22x1_ASAP7_75t_R ALU___U291 ( .A1(ALU__N172), .A2(ALU__n1564), .B1(ALU__N281), .B2(ALU__n1535), .Y(
        n192) );
  BUFx12f_ASAP7_75t_R ALU___U293 ( .A(ALU__n390), .Y(ALU__n348) );
  BUFx12f_ASAP7_75t_R ALU___U297 ( .A(ALU__n659), .Y(ALU__n349) );
  BUFx12f_ASAP7_75t_R ALU___U298 ( .A(ALU__n377), .Y(ALU__n350) );
  BUFx12f_ASAP7_75t_R ALU___U300 ( .A(ALU__n377), .Y(ALU__n351) );
  BUFx16f_ASAP7_75t_R ALU___U304 ( .A(ALU__n1175), .Y(ALU__n352) );
  CKINVDCx10_ASAP7_75t_R ALU___U305 ( .A(ALU__n352), .Y(ALU__n1482) );
  BUFx16f_ASAP7_75t_R ALU___U307 ( .A(ALU__n675), .Y(ALU__n353) );
  CKINVDCx10_ASAP7_75t_R ALU___U311 ( .A(ALU__n353), .Y(ALU__n1622) );
  BUFx12f_ASAP7_75t_R ALU___U312 ( .A(ALU__n1295), .Y(ALU__n675) );
  BUFx3_ASAP7_75t_R ALU___U314 ( .A(ALU__n355), .Y(ALU__n354) );
  BUFx2_ASAP7_75t_R ALU___U318 ( .A(ALU__n270), .Y(ALU__n355) );
  BUFx4f_ASAP7_75t_R ALU___U319 ( .A(ALU__n354), .Y(ALU__n638) );
  BUFx4f_ASAP7_75t_R ALU___U321 ( .A(ALU__n357), .Y(ALU__n356) );
  BUFx3_ASAP7_75t_R ALU___U325 ( .A(ALU__n10), .Y(ALU__n357) );
  BUFx2_ASAP7_75t_R ALU___U326 ( .A(ALU__n381), .Y(ALU__n358) );
  BUFx4f_ASAP7_75t_R ALU___U328 ( .A(ALU__n360), .Y(ALU__n359) );
  INVx2_ASAP7_75t_R ALU___U332 ( .A(ALU__n359), .Y(ALU__n1003) );
  BUFx12f_ASAP7_75t_R ALU___U333 ( .A(ALU__n686), .Y(ALU__n361) );
  BUFx12f_ASAP7_75t_R ALU___U335 ( .A(ALU__n686), .Y(ALU__n362) );
  INVx6_ASAP7_75t_R ALU___U339 ( .A(ALU__n845), .Y(ALU__n1392) );
  INVx6_ASAP7_75t_R ALU___U340 ( .A(ALU__n1320), .Y(ALU__n1390) );
  BUFx2_ASAP7_75t_R ALU___U342 ( .A(ALU__n300), .Y(ALU__n363) );
  BUFx2_ASAP7_75t_R ALU___U345 ( .A(ALU__n312), .Y(ALU__n364) );
  BUFx2_ASAP7_75t_R ALU___U347 ( .A(ALU__n152), .Y(ALU__n365) );
  BUFx2_ASAP7_75t_R ALU___U352 ( .A(ALU__n308), .Y(ALU__n366) );
  BUFx12f_ASAP7_75t_R ALU___U353 ( .A(n341), .Y(ALU__n367) );
  BUFx12f_ASAP7_75t_R ALU___U354 ( .A(n341), .Y(ALU__n368) );
  BUFx3_ASAP7_75t_R ALU___U356 ( .A(ALU__n370), .Y(ALU__n369) );
  BUFx2_ASAP7_75t_R ALU___U357 ( .A(ALU__n161), .Y(ALU__n370) );
  BUFx3_ASAP7_75t_R ALU___U358 ( .A(ALU__n372), .Y(ALU__n371) );
  BUFx2_ASAP7_75t_R ALU___U359 ( .A(ALU__n159), .Y(ALU__n372) );
  BUFx4f_ASAP7_75t_R ALU___U360 ( .A(ALU__n374), .Y(ALU__n373) );
  INVx2_ASAP7_75t_R ALU___U361 ( .A(ALU__n373), .Y(ALU__n937) );
  BUFx12f_ASAP7_75t_R ALU___U362 ( .A(ALU__n1327), .Y(ALU__n375) );
  BUFx12f_ASAP7_75t_R ALU___U363 ( .A(ALU__n1327), .Y(ALU__n376) );
  BUFx12f_ASAP7_75t_R ALU___U364 ( .A(ALU__n649), .Y(ALU__n377) );
  CKINVDCx10_ASAP7_75t_R ALU___U365 ( .A(ALU__n676), .Y(ALU__n1621) );
  BUFx12f_ASAP7_75t_R ALU___U366 ( .A(ALU__n379), .Y(ALU__n378) );
  BUFx12f_ASAP7_75t_R ALU___U367 ( .A(ALU__n1617), .Y(ALU__n379) );
  OR2x2_ASAP7_75t_R ALU___U368 ( .A(ALU__n358), .B(ALU__n1427), .Y(ALU__n380) );
  OR2x2_ASAP7_75t_R ALU___U369 ( .A(ALU_ctl[3]), .B(ALU__n646), .Y(ALU__n381) );
  BUFx2_ASAP7_75t_R ALU___U370 ( .A(ALU__n1428), .Y(ALU__n382) );
  INVx6_ASAP7_75t_R ALU___U371 ( .A(ALU__n378), .Y(ALU__n1426) );
  INVx1_ASAP7_75t_R ALU___U372 ( .A(ALU__n382), .Y(ALU__n1427) );
  CKINVDCx14_ASAP7_75t_R ALU___U373 ( .A(ALU__n396), .Y(ALU__n394) );
  BUFx4f_ASAP7_75t_R ALU___U374 ( .A(ALU__n384), .Y(ALU__n383) );
  BUFx3_ASAP7_75t_R ALU___U375 ( .A(ALU__n90), .Y(ALU__n384) );
  AO22x1_ASAP7_75t_R ALU___U376 ( .A1(ALU__N168), .A2(ALU__n1556), .B1(ALU__N277), .B2(ALU__n1533), .Y(
        n216) );
  BUFx2_ASAP7_75t_R ALU___U377 ( .A(ALU__n1651), .Y(ALU__n385) );
  BUFx3_ASAP7_75t_R ALU___U378 ( .A(ALU__n387), .Y(ALU__n386) );
  BUFx2_ASAP7_75t_R ALU___U379 ( .A(ALU__n1650), .Y(ALU__n387) );
  BUFx3_ASAP7_75t_R ALU___U380 ( .A(ALU__n389), .Y(ALU__n388) );
  BUFx2_ASAP7_75t_R ALU___U381 ( .A(ALU__n1652), .Y(ALU__n389) );
  AO221x1_ASAP7_75t_R ALU___U382 ( .A1(n1174), .A2(ALU__n1747), .B1(
        n1060), .B2(ALU__n1746), .C(ALU__n737), .Y(ALU__n1650) );
  AO221x1_ASAP7_75t_R ALU___U383 ( .A1(n973), .A2(ALU__n1194), .B1(
        n1233), .B2(ALU__n1682), .C(ALU__n385), .Y(ALU__n1652) );
  BUFx12f_ASAP7_75t_R ALU___U384 ( .A(ALU__n781), .Y(ALU__n390) );
  BUFx12f_ASAP7_75t_R ALU___U385 ( .A(ALU__n1067), .Y(ALU__n391) );
  BUFx3_ASAP7_75t_R ALU___U386 ( .A(ALU__n393), .Y(ALU__n392) );
  BUFx2_ASAP7_75t_R ALU___U387 ( .A(ALU__n252), .Y(ALU__n393) );
  AO22x2_ASAP7_75t_R ALU___U388 ( .A1(ALU__N162), .A2(ALU__n1560), .B1(ALU__N271), .B2(ALU__n1530), .Y(
        n252) );
  BUFx4f_ASAP7_75t_R ALU___U389 ( .A(ALU__n392), .Y(ALU__n534) );
  CKINVDCx14_ASAP7_75t_R ALU___U390 ( .A(ALU__n701), .Y(ALU__n1518) );
  CKINVDCx16_ASAP7_75t_R ALU___U391 ( .A(ALU__n394), .Y(ALU__n395) );
  BUFx16f_ASAP7_75t_R ALU___U392 ( .A(ALU__n1338), .Y(ALU__n396) );
  CKINVDCx16_ASAP7_75t_R ALU___U393 ( .A(ALU__n395), .Y(ALU__n1481) );
  BUFx12f_ASAP7_75t_R ALU___U394 ( .A(ALU__n41), .Y(ALU__n1338) );
  BUFx16f_ASAP7_75t_R ALU___U395 ( .A(ALU__n1365), .Y(ALU__n397) );
  CKINVDCx16_ASAP7_75t_R ALU___U396 ( .A(ALU__n397), .Y(ALU__n1619) );
  BUFx12f_ASAP7_75t_R ALU___U397 ( .A(ALU__n1294), .Y(ALU__n1365) );
  BUFx12f_ASAP7_75t_R ALU___U398 ( .A(ALU__n54), .Y(ALU__n398) );
  BUFx12f_ASAP7_75t_R ALU___U399 ( .A(ALU__n54), .Y(ALU__n399) );
  BUFx12f_ASAP7_75t_R ALU___U400 ( .A(ALU__n857), .Y(ALU__n400) );
  INVx5_ASAP7_75t_R ALU___U401 ( .A(ALU__n399), .Y(ALU__n1593) );
  BUFx12f_ASAP7_75t_R ALU___U402 ( .A(ALU__n859), .Y(ALU__n857) );
  BUFx3_ASAP7_75t_R ALU___U403 ( .A(ALU__n402), .Y(ALU__n401) );
  BUFx2_ASAP7_75t_R ALU___U404 ( .A(ALU__n204), .Y(ALU__n402) );
  BUFx4f_ASAP7_75t_R ALU___U405 ( .A(ALU__n401), .Y(ALU__n541) );
  BUFx4f_ASAP7_75t_R ALU___U406 ( .A(ALU__n404), .Y(ALU__n403) );
  BUFx3_ASAP7_75t_R ALU___U407 ( .A(ALU__n74), .Y(ALU__n404) );
  BUFx2_ASAP7_75t_R ALU___U408 ( .A(ALU__n1655), .Y(ALU__n405) );
  BUFx2_ASAP7_75t_R ALU___U409 ( .A(ALU__n1653), .Y(ALU__n406) );
  BUFx3_ASAP7_75t_R ALU___U410 ( .A(ALU__n408), .Y(ALU__n407) );
  BUFx2_ASAP7_75t_R ALU___U411 ( .A(ALU__n1654), .Y(ALU__n408) );
  AO221x1_ASAP7_75t_R ALU___U412 ( .A1(n929), .A2(ALU__n1680), .B1(
        n1114), .B2(ALU__n1235), .C(ALU__n406), .Y(ALU__n1654) );
  BUFx12f_ASAP7_75t_R ALU___U413 ( .A(n435), .Y(ALU__n409) );
  BUFx12f_ASAP7_75t_R ALU___U414 ( .A(n435), .Y(ALU__n410) );
  CKINVDCx14_ASAP7_75t_R ALU___U415 ( .A(ALU__n420), .Y(ALU__n418) );
  BUFx3_ASAP7_75t_R ALU___U416 ( .A(ALU__n412), .Y(ALU__n411) );
  BUFx2_ASAP7_75t_R ALU___U417 ( .A(ALU__n197), .Y(ALU__n412) );
  BUFx3_ASAP7_75t_R ALU___U418 ( .A(ALU__n414), .Y(ALU__n413) );
  BUFx2_ASAP7_75t_R ALU___U419 ( .A(ALU__n195), .Y(ALU__n414) );
  BUFx12f_ASAP7_75t_R ALU___U420 ( .A(ALU__n1578), .Y(ALU__n1379) );
  BUFx12f_ASAP7_75t_R ALU___U421 ( .A(ALU__n807), .Y(ALU__n1578) );
  INVx4_ASAP7_75t_R ALU___U422 ( .A(ALU__n1571), .Y(ALU__n1566) );
  INVx4_ASAP7_75t_R ALU___U423 ( .A(ALU__n1572), .Y(ALU__n1565) );
  BUFx6f_ASAP7_75t_R ALU___U424 ( .A(ALU__n66), .Y(ALU__n415) );
  BUFx3_ASAP7_75t_R ALU___U425 ( .A(ALU__n133), .Y(ALU__n416) );
  OR4x1_ASAP7_75t_R ALU___U426 ( .A(ALU__n1349), .B(ALU__n1406), .C(ALU_ctl[3]), .D(
        ALU_ctl[1]), .Y(ALU__n133) );
  BUFx12f_ASAP7_75t_R ALU___U427 ( .A(ALU__n415), .Y(ALU__n808) );
  CKINVDCx16_ASAP7_75t_R ALU___U428 ( .A(ALU__n418), .Y(ALU__n419) );
  BUFx16f_ASAP7_75t_R ALU___U429 ( .A(ALU__n1340), .Y(ALU__n420) );
  CKINVDCx16_ASAP7_75t_R ALU___U430 ( .A(ALU__n419), .Y(ALU__n1484) );
  BUFx12f_ASAP7_75t_R ALU___U431 ( .A(ALU__n1055), .Y(ALU__n1340) );
  BUFx3_ASAP7_75t_R ALU___U432 ( .A(ALU__n422), .Y(ALU__n421) );
  BUFx2_ASAP7_75t_R ALU___U433 ( .A(ALU__n167), .Y(ALU__n422) );
  BUFx3_ASAP7_75t_R ALU___U434 ( .A(ALU__n424), .Y(ALU__n423) );
  BUFx2_ASAP7_75t_R ALU___U435 ( .A(ALU__n165), .Y(ALU__n424) );
  BUFx2_ASAP7_75t_R ALU___U436 ( .A(ALU__n1667), .Y(ALU__n425) );
  BUFx2_ASAP7_75t_R ALU___U437 ( .A(ALU__n1665), .Y(ALU__n426) );
  BUFx3_ASAP7_75t_R ALU___U438 ( .A(ALU__n428), .Y(ALU__n427) );
  BUFx2_ASAP7_75t_R ALU___U439 ( .A(ALU__n1666), .Y(ALU__n428) );
  AO221x1_ASAP7_75t_R ALU___U440 ( .A1(n1068), .A2(ALU__n1690), .B1(ALU__n1037), 
        .B2(ALU__n1298), .C(ALU__n426), .Y(ALU__n1666) );
  INVx3_ASAP7_75t_R ALU___U441 ( .A(ALU__n1539), .Y(ALU__n1538) );
  INVx4_ASAP7_75t_R ALU___U442 ( .A(ALU__n1543), .Y(ALU__n1533) );
  BUFx6f_ASAP7_75t_R ALU___U443 ( .A(ALU__n67), .Y(ALU__n429) );
  BUFx3_ASAP7_75t_R ALU___U444 ( .A(ALU__n132), .Y(ALU__n430) );
  OR4x1_ASAP7_75t_R ALU___U445 ( .A(ALU__n1349), .B(ALU__n988), .C(ALU_ctl[3]), .D(ALU__n646), 
        .Y(ALU__n132) );
  BUFx12f_ASAP7_75t_R ALU___U446 ( .A(ALU__n429), .Y(ALU__n854) );
  BUFx12f_ASAP7_75t_R ALU___U447 ( .A(ALU__n687), .Y(ALU__n432) );
  BUFx2_ASAP7_75t_R ALU___U448 ( .A(ALU__n266), .Y(ALU__n433) );
  BUFx3_ASAP7_75t_R ALU___U449 ( .A(ALU__n435), .Y(ALU__n434) );
  BUFx2_ASAP7_75t_R ALU___U450 ( .A(ALU__n191), .Y(ALU__n435) );
  BUFx3_ASAP7_75t_R ALU___U451 ( .A(ALU__n437), .Y(ALU__n436) );
  BUFx2_ASAP7_75t_R ALU___U452 ( .A(ALU__n189), .Y(ALU__n437) );
  BUFx3_ASAP7_75t_R ALU___U453 ( .A(ALU__n439), .Y(ALU__n438) );
  BUFx2_ASAP7_75t_R ALU___U454 ( .A(ALU__n275), .Y(ALU__n439) );
  BUFx3_ASAP7_75t_R ALU___U455 ( .A(ALU__n441), .Y(ALU__n440) );
  BUFx2_ASAP7_75t_R ALU___U456 ( .A(ALU__n273), .Y(ALU__n441) );
  BUFx12f_ASAP7_75t_R ALU___U457 ( .A(ALU__n1379), .Y(ALU__n1581) );
  INVx4_ASAP7_75t_R ALU___U458 ( .A(ALU__n1574), .Y(ALU__n1563) );
  INVx3_ASAP7_75t_R ALU___U459 ( .A(ALU__n1569), .Y(ALU__n1568) );
  INVx2_ASAP7_75t_R ALU___U460 ( .A(ALU__n1551), .Y(ALU__n1526) );
  BUFx12f_ASAP7_75t_R ALU___U461 ( .A(ALU__n1356), .Y(ALU__n1551) );
  BUFx2_ASAP7_75t_R ALU___U462 ( .A(ALU__n146), .Y(ALU__n442) );
  BUFx2_ASAP7_75t_R ALU___U463 ( .A(ALU__n306), .Y(ALU__n443) );
  INVx5_ASAP7_75t_R ALU___U464 ( .A(ALU__n708), .Y(ALU__n1386) );
  BUFx3_ASAP7_75t_R ALU___U465 ( .A(ALU__n445), .Y(ALU__n444) );
  BUFx2_ASAP7_75t_R ALU___U466 ( .A(ALU__n185), .Y(ALU__n445) );
  BUFx3_ASAP7_75t_R ALU___U467 ( .A(ALU__n447), .Y(ALU__n446) );
  BUFx2_ASAP7_75t_R ALU___U468 ( .A(ALU__n183), .Y(ALU__n447) );
  AO22x2_ASAP7_75t_R ALU___U469 ( .A1(ALU__N314), .A2(ALU__n1518), .B1(ALU__N346), .B2(ALU__n1505), .Y(
        n184) );
  BUFx3_ASAP7_75t_R ALU___U470 ( .A(ALU__n449), .Y(ALU__n448) );
  BUFx2_ASAP7_75t_R ALU___U471 ( .A(ALU__n215), .Y(ALU__n449) );
  BUFx3_ASAP7_75t_R ALU___U472 ( .A(ALU__n451), .Y(ALU__n450) );
  BUFx2_ASAP7_75t_R ALU___U473 ( .A(ALU__n213), .Y(ALU__n451) );
  BUFx3_ASAP7_75t_R ALU___U474 ( .A(ALU__n453), .Y(ALU__n452) );
  BUFx2_ASAP7_75t_R ALU___U475 ( .A(ALU__n281), .Y(ALU__n453) );
  BUFx3_ASAP7_75t_R ALU___U476 ( .A(ALU__n455), .Y(ALU__n454) );
  BUFx2_ASAP7_75t_R ALU___U477 ( .A(ALU__n279), .Y(ALU__n455) );
  BUFx4f_ASAP7_75t_R ALU___U478 ( .A(ALU__n457), .Y(ALU__n456) );
  BUFx3_ASAP7_75t_R ALU___U479 ( .A(ALU__n76), .Y(ALU__n457) );
  INVx4_ASAP7_75t_R ALU___U480 ( .A(n701), .Y(ALU__n1690) );
  BUFx2_ASAP7_75t_R ALU___U481 ( .A(ALU__n135), .Y(ALU__n458) );
  BUFx12f_ASAP7_75t_R ALU___U482 ( .A(ALU__n460), .Y(ALU__n459) );
  BUFx12f_ASAP7_75t_R ALU___U483 ( .A(ALU__n1513), .Y(ALU__n460) );
  INVx6_ASAP7_75t_R ALU___U484 ( .A(ALU__n459), .Y(ALU__n1342) );
  BUFx12f_ASAP7_75t_R ALU___U485 ( .A(ALU__n463), .Y(ALU__n461) );
  BUFx12f_ASAP7_75t_R ALU___U486 ( .A(ALU__n463), .Y(ALU__n462) );
  BUFx12f_ASAP7_75t_R ALU___U487 ( .A(ALU__n762), .Y(ALU__n463) );
  BUFx16f_ASAP7_75t_R ALU___U488 ( .A(ALU__n498), .Y(ALU__n464) );
  BUFx12f_ASAP7_75t_R ALU___U489 ( .A(ALU__n703), .Y(ALU__n498) );
  CKINVDCx14_ASAP7_75t_R ALU___U490 ( .A(ALU__n496), .Y(ALU__n494) );
  BUFx12f_ASAP7_75t_R ALU___U491 ( .A(ALU__n50), .Y(ALU__n465) );
  BUFx12f_ASAP7_75t_R ALU___U492 ( .A(ALU__n44), .Y(ALU__n466) );
  BUFx12f_ASAP7_75t_R ALU___U493 ( .A(ALU__n745), .Y(ALU__n467) );
  CKINVDCx5p33_ASAP7_75t_R ALU___U494 ( .A(ALU__n466), .Y(ALU__n1605) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U495 ( .A(ALU__n465), .Y(ALU__n1603) );
  BUFx12f_ASAP7_75t_R ALU___U496 ( .A(ALU__n343), .Y(ALU__n745) );
  INVx2_ASAP7_75t_R ALU___U497 ( .A(ALU__n1550), .Y(ALU__n1527) );
  BUFx12f_ASAP7_75t_R ALU___U498 ( .A(ALU__n1551), .Y(ALU__n1550) );
  BUFx12f_ASAP7_75t_R ALU___U499 ( .A(ALU__n9), .Y(ALU__n1576) );
  BUFx4f_ASAP7_75t_R ALU___U500 ( .A(ALU__n9), .Y(ALU__n1579) );
  BUFx3_ASAP7_75t_R ALU___U501 ( .A(ALU__n470), .Y(ALU__n469) );
  BUFx2_ASAP7_75t_R ALU___U502 ( .A(ALU__n137), .Y(ALU__n470) );
  BUFx2_ASAP7_75t_R ALU___U503 ( .A(ALU__n1407), .Y(ALU__n471) );
  BUFx2_ASAP7_75t_R ALU___U504 ( .A(ALU__n1408), .Y(ALU__n472) );
  INVx6_ASAP7_75t_R ALU___U505 ( .A(ALU__n1072), .Y(ALU__n1420) );
  INVx6_ASAP7_75t_R ALU___U506 ( .A(ALU__n1376), .Y(ALU__n1415) );
  BUFx2_ASAP7_75t_R ALU___U507 ( .A(ALU__n194), .Y(ALU__n473) );
  BUFx2_ASAP7_75t_R ALU___U508 ( .A(ALU__N356), .Y(ALU__n474) );
  BUFx2_ASAP7_75t_R ALU___U509 ( .A(ALU__n1170), .Y(ALU__n475) );
  BUFx3_ASAP7_75t_R ALU___U510 ( .A(ALU__n477), .Y(ALU__n476) );
  BUFx2_ASAP7_75t_R ALU___U511 ( .A(ALU__n321), .Y(ALU__n477) );
  AND3x1_ASAP7_75t_R ALU___U512 ( .A(ALU__n1172), .B(ALU__n1173), .C(ALU__n1171), .Y(ALU__N356) );
  INVx6_ASAP7_75t_R ALU___U513 ( .A(ALU__n485), .Y(ALU__n1744) );
  INVx5_ASAP7_75t_R ALU___U514 ( .A(ALU__n838), .Y(ALU__n1358) );
  BUFx3_ASAP7_75t_R ALU___U515 ( .A(ALU__n479), .Y(ALU__n478) );
  BUFx2_ASAP7_75t_R ALU___U516 ( .A(ALU__n299), .Y(ALU__n479) );
  BUFx3_ASAP7_75t_R ALU___U517 ( .A(ALU__n481), .Y(ALU__n480) );
  BUFx2_ASAP7_75t_R ALU___U518 ( .A(ALU__n297), .Y(ALU__n481) );
  BUFx2_ASAP7_75t_R ALU___U519 ( .A(ALU__n307), .Y(ALU__n482) );
  INVx5_ASAP7_75t_R ALU___U520 ( .A(ALU__n1199), .Y(ALU__n1421) );
  CKINVDCx10_ASAP7_75t_R ALU___U521 ( .A(ALU__n1535), .Y(ALU__n483) );
  BUFx12f_ASAP7_75t_R ALU___U522 ( .A(ALU__n483), .Y(ALU__n1545) );
  BUFx4f_ASAP7_75t_R ALU___U523 ( .A(ALU__n483), .Y(ALU__n1548) );
  BUFx16f_ASAP7_75t_R ALU___U524 ( .A(ALU__n1167), .Y(ALU__n1356) );
  INVx2_ASAP7_75t_R ALU___U525 ( .A(ALU__n1579), .Y(ALU__n1559) );
  BUFx2_ASAP7_75t_R ALU___U526 ( .A(ALU__n1743), .Y(ALU__n484) );
  BUFx12f_ASAP7_75t_R ALU___U527 ( .A(ALU__n683), .Y(ALU__n485) );
  BUFx12f_ASAP7_75t_R ALU___U528 ( .A(ALU__n488), .Y(ALU__n486) );
  BUFx12f_ASAP7_75t_R ALU___U529 ( .A(ALU__n489), .Y(ALU__n487) );
  BUFx12f_ASAP7_75t_R ALU___U530 ( .A(ALU__n574), .Y(ALU__n488) );
  BUFx12f_ASAP7_75t_R ALU___U531 ( .A(ALU__n574), .Y(ALU__n489) );
  BUFx3_ASAP7_75t_R ALU___U532 ( .A(ALU__n613), .Y(ALU__n490) );
  CKINVDCx10_ASAP7_75t_R ALU___U533 ( .A(ALU__n614), .Y(ALU__n1018) );
  INVx6_ASAP7_75t_R ALU___U534 ( .A(ALU__n609), .Y(ALU__n981) );
  BUFx3_ASAP7_75t_R ALU___U535 ( .A(ALU__n492), .Y(ALU__n491) );
  BUFx2_ASAP7_75t_R ALU___U536 ( .A(ALU__n276), .Y(ALU__n492) );
  AO22x2_ASAP7_75t_R ALU___U537 ( .A1(ALU__N158), .A2(ALU__n1559), .B1(ALU__N267), .B2(ALU__n1529), .Y(
        n276) );
  BUFx4f_ASAP7_75t_R ALU___U538 ( .A(ALU__n491), .Y(ALU__n729) );
  BUFx2_ASAP7_75t_R ALU___U539 ( .A(ALU__n330), .Y(ALU__n493) );
  AND3x1_ASAP7_75t_R ALU___U540 ( .A(ALU_ctl[1]), .B(ALU_ctl[0]), .C(ALU__n646), 
        .Y(ALU__n330) );
  CKINVDCx16_ASAP7_75t_R ALU___U541 ( .A(ALU__n494), .Y(ALU__n495) );
  BUFx16f_ASAP7_75t_R ALU___U542 ( .A(ALU__n1341), .Y(ALU__n496) );
  CKINVDCx16_ASAP7_75t_R ALU___U543 ( .A(ALU__n495), .Y(ALU__n1485) );
  BUFx12f_ASAP7_75t_R ALU___U544 ( .A(ALU__n1493), .Y(ALU__n1341) );
  BUFx16f_ASAP7_75t_R ALU___U545 ( .A(ALU__n647), .Y(ALU__n497) );
  INVx13_ASAP7_75t_R ALU___U546 ( .A(ALU__n497), .Y(ALU__n1517) );
  BUFx12f_ASAP7_75t_R ALU___U547 ( .A(ALU__n350), .Y(ALU__n647) );
  BUFx12f_ASAP7_75t_R ALU___U548 ( .A(ALU__n1627), .Y(ALU__n703) );
  BUFx12f_ASAP7_75t_R ALU___U549 ( .A(ALU__n22), .Y(ALU__n499) );
  BUFx12f_ASAP7_75t_R ALU___U550 ( .A(ALU__n23), .Y(ALU__n500) );
  BUFx12f_ASAP7_75t_R ALU___U551 ( .A(ALU__n106), .Y(ALU__n1610) );
  BUFx12f_ASAP7_75t_R ALU___U552 ( .A(ALU__n1615), .Y(ALU__n1613) );
  BUFx12f_ASAP7_75t_R ALU___U553 ( .A(ALU__n1616), .Y(ALU__n1606) );
  BUFx3_ASAP7_75t_R ALU___U554 ( .A(ALU__n502), .Y(ALU__n501) );
  BUFx2_ASAP7_75t_R ALU___U555 ( .A(ALU__n144), .Y(ALU__n502) );
  BUFx4f_ASAP7_75t_R ALU___U556 ( .A(ALU__n501), .Y(ALU__n525) );
  BUFx12f_ASAP7_75t_R ALU___U557 ( .A(ALU__n782), .Y(ALU__n503) );
  BUFx6f_ASAP7_75t_R ALU___U558 ( .A(ALU__n971), .Y(ALU__n504) );
  BUFx12f_ASAP7_75t_R ALU___U559 ( .A(ALU__n971), .Y(ALU__n505) );
  BUFx3_ASAP7_75t_R ALU___U560 ( .A(ALU__n507), .Y(ALU__n506) );
  BUFx2_ASAP7_75t_R ALU___U561 ( .A(ALU__n1677), .Y(ALU__n507) );
  BUFx2_ASAP7_75t_R ALU___U562 ( .A(ALU__n272), .Y(ALU__n508) );
  BUFx2_ASAP7_75t_R ALU___U563 ( .A(ALU__n318), .Y(ALU__n509) );
  BUFx3_ASAP7_75t_R ALU___U564 ( .A(ALU__n511), .Y(ALU__n510) );
  BUFx2_ASAP7_75t_R ALU___U565 ( .A(ALU__n282), .Y(ALU__n511) );
  AO22x2_ASAP7_75t_R ALU___U566 ( .A1(ALU__N157), .A2(ALU__n1558), .B1(ALU__N266), .B2(ALU__n1528), .Y(
        n282) );
  BUFx4f_ASAP7_75t_R ALU___U567 ( .A(ALU__n510), .Y(ALU__n821) );
  BUFx2_ASAP7_75t_R ALU___U568 ( .A(ALU__n182), .Y(ALU__n512) );
  BUFx2_ASAP7_75t_R ALU___U569 ( .A(ALU__n514), .Y(ALU__n513) );
  BUFx2_ASAP7_75t_R ALU___U570 ( .A(ALU__n206), .Y(ALU__n514) );
  BUFx2_ASAP7_75t_R ALU___U571 ( .A(ALU__n242), .Y(ALU__n515) );
  BUFx2_ASAP7_75t_R ALU___U572 ( .A(ALU__n254), .Y(ALU__n516) );
  BUFx4f_ASAP7_75t_R ALU___U573 ( .A(ALU__n518), .Y(ALU__n517) );
  BUFx3_ASAP7_75t_R ALU___U574 ( .A(ALU__n364), .Y(ALU__n518) );
  BUFx2_ASAP7_75t_R ALU___U575 ( .A(ALU__n199), .Y(ALU__n519) );
  INVx6_ASAP7_75t_R ALU___U576 ( .A(ALU__n1764), .Y(ALU__n1335) );
  BUFx3_ASAP7_75t_R ALU___U577 ( .A(ALU__n521), .Y(ALU__n520) );
  BUFx2_ASAP7_75t_R ALU___U578 ( .A(ALU__n128), .Y(ALU__n521) );
  BUFx3_ASAP7_75t_R ALU___U579 ( .A(ALU__n523), .Y(ALU__n522) );
  BUFx2_ASAP7_75t_R ALU___U580 ( .A(ALU__n126), .Y(ALU__n523) );
  INVx6_ASAP7_75t_R ALU___U581 ( .A(ALU__n1736), .Y(ALU__n1349) );
  BUFx12f_ASAP7_75t_R ALU___U582 ( .A(ALU_ctl[0]), .Y(ALU__n1736) );
  BUFx4f_ASAP7_75t_R ALU___U583 ( .A(ALU__n525), .Y(ALU__n524) );
  INVx2_ASAP7_75t_R ALU___U584 ( .A(ALU__n524), .Y(ALU__n1063) );
  BUFx3_ASAP7_75t_R ALU___U585 ( .A(ALU__n544), .Y(ALU__n526) );
  INVx6_ASAP7_75t_R ALU___U586 ( .A(ALU__n1768), .Y(ALU__n1385) );
  INVx6_ASAP7_75t_R ALU___U587 ( .A(ALU__n724), .Y(ALU__n1387) );
  BUFx4f_ASAP7_75t_R ALU___U588 ( .A(ALU__n528), .Y(ALU__n527) );
  BUFx3_ASAP7_75t_R ALU___U589 ( .A(ALU__n324), .Y(ALU__n528) );
  BUFx2_ASAP7_75t_R ALU___U590 ( .A(ALU__n1422), .Y(ALU__n1024) );
  INVx1_ASAP7_75t_R ALU___U591 ( .A(ALU__n1024), .Y(ALU__n529) );
  BUFx2_ASAP7_75t_R ALU___U592 ( .A(ALU__n164), .Y(ALU__n530) );
  BUFx2_ASAP7_75t_R ALU___U593 ( .A(ALU__n218), .Y(ALU__n531) );
  BUFx2_ASAP7_75t_R ALU___U594 ( .A(ALU__n508), .Y(ALU__n532) );
  BUFx4f_ASAP7_75t_R ALU___U595 ( .A(ALU__n534), .Y(ALU__n533) );
  INVx2_ASAP7_75t_R ALU___U596 ( .A(ALU__n533), .Y(ALU__n1409) );
  BUFx3_ASAP7_75t_R ALU___U597 ( .A(ALU__n536), .Y(ALU__n535) );
  BUFx2_ASAP7_75t_R ALU___U598 ( .A(ALU__n227), .Y(ALU__n536) );
  BUFx3_ASAP7_75t_R ALU___U599 ( .A(ALU__n538), .Y(ALU__n537) );
  BUFx2_ASAP7_75t_R ALU___U600 ( .A(ALU__n225), .Y(ALU__n538) );
  BUFx2_ASAP7_75t_R ALU___U601 ( .A(ALU__n150), .Y(ALU__n539) );
  BUFx4f_ASAP7_75t_R ALU___U602 ( .A(ALU__n541), .Y(ALU__n540) );
  INVx2_ASAP7_75t_R ALU___U603 ( .A(ALU__n540), .Y(ALU__n1234) );
  BUFx12f_ASAP7_75t_R ALU___U604 ( .A(ALU__n543), .Y(ALU__n542) );
  BUFx12f_ASAP7_75t_R ALU___U605 ( .A(ALU__n575), .Y(ALU__n543) );
  INVx6_ASAP7_75t_R ALU___U606 ( .A(ALU__n748), .Y(ALU__n1359) );
  BUFx2_ASAP7_75t_R ALU___U607 ( .A(ALU__n288), .Y(ALU__n544) );
  AO22x2_ASAP7_75t_R ALU___U608 ( .A1(ALU__N156), .A2(ALU__n1558), .B1(ALU__N265), .B2(ALU__n1528), .Y(
        n288) );
  INVx2_ASAP7_75t_R ALU___U609 ( .A(ALU__n1108), .Y(ALU__n1132) );
  BUFx4f_ASAP7_75t_R ALU___U610 ( .A(ALU__n526), .Y(ALU__n1108) );
  BUFx2_ASAP7_75t_R ALU___U611 ( .A(ALU__n546), .Y(ALU__n545) );
  BUFx2_ASAP7_75t_R ALU___U612 ( .A(ALU__n278), .Y(ALU__n546) );
  BUFx4f_ASAP7_75t_R ALU___U613 ( .A(ALU__n548), .Y(ALU__n547) );
  BUFx3_ASAP7_75t_R ALU___U614 ( .A(ALU__n363), .Y(ALU__n548) );
  BUFx4f_ASAP7_75t_R ALU___U615 ( .A(ALU__n550), .Y(ALU__n549) );
  BUFx3_ASAP7_75t_R ALU___U616 ( .A(ALU__n509), .Y(ALU__n550) );
  BUFx3_ASAP7_75t_R ALU___U617 ( .A(ALU__n552), .Y(ALU__n551) );
  BUFx2_ASAP7_75t_R ALU___U618 ( .A(ALU__n155), .Y(ALU__n552) );
  BUFx3_ASAP7_75t_R ALU___U619 ( .A(ALU__n554), .Y(ALU__n553) );
  BUFx2_ASAP7_75t_R ALU___U620 ( .A(ALU__n153), .Y(ALU__n554) );
  BUFx3_ASAP7_75t_R ALU___U621 ( .A(ALU__n556), .Y(ALU__n555) );
  BUFx2_ASAP7_75t_R ALU___U622 ( .A(ALU__n209), .Y(ALU__n556) );
  BUFx3_ASAP7_75t_R ALU___U623 ( .A(ALU__n558), .Y(ALU__n557) );
  BUFx2_ASAP7_75t_R ALU___U624 ( .A(ALU__n207), .Y(ALU__n558) );
  BUFx3_ASAP7_75t_R ALU___U625 ( .A(ALU__n560), .Y(ALU__n559) );
  BUFx2_ASAP7_75t_R ALU___U626 ( .A(ALU__n305), .Y(ALU__n560) );
  BUFx3_ASAP7_75t_R ALU___U627 ( .A(ALU__n562), .Y(ALU__n561) );
  BUFx2_ASAP7_75t_R ALU___U628 ( .A(ALU__n303), .Y(ALU__n562) );
  BUFx2_ASAP7_75t_R ALU___U629 ( .A(ALU__n181), .Y(ALU__n563) );
  BUFx2_ASAP7_75t_R ALU___U630 ( .A(ALU__n241), .Y(ALU__n564) );
  INVx5_ASAP7_75t_R ALU___U631 ( .A(ALU__n1237), .Y(ALU__n1337) );
  BUFx4f_ASAP7_75t_R ALU___U632 ( .A(ALU__n566), .Y(ALU__n565) );
  BUFx3_ASAP7_75t_R ALU___U633 ( .A(ALU__n539), .Y(ALU__n566) );
  BUFx2_ASAP7_75t_R ALU___U634 ( .A(ALU__n131), .Y(ALU__n567) );
  AO22x2_ASAP7_75t_R ALU___U635 ( .A1(ALU__N181), .A2(ALU__n1568), .B1(ALU__N290), .B2(ALU__n1538), .Y(
        n131) );
  AO22x2_ASAP7_75t_R ALU___U636 ( .A1(ALU__N175), .A2(ALU__n1565), .B1(ALU__N284), .B2(ALU__n1536), .Y(
        n174) );
  INVx2_ASAP7_75t_R ALU___U637 ( .A(ALU__n344), .Y(ALU__n568) );
  BUFx2_ASAP7_75t_R ALU___U638 ( .A(ALU__n234), .Y(ALU__n662) );
  INVx1_ASAP7_75t_R ALU___U639 ( .A(ALU__n662), .Y(ALU__n569) );
  BUFx12f_ASAP7_75t_R ALU___U640 ( .A(ALU__n571), .Y(ALU__n570) );
  BUFx12f_ASAP7_75t_R ALU___U641 ( .A(ALU__n1777), .Y(ALU__n571) );
  INVx6_ASAP7_75t_R ALU___U642 ( .A(ALU__n1039), .Y(ALU__n1360) );
  BUFx12f_ASAP7_75t_R ALU___U643 ( .A(ALU__n658), .Y(ALU__n572) );
  BUFx12f_ASAP7_75t_R ALU___U644 ( .A(ALU__n487), .Y(ALU__n573) );
  BUFx12f_ASAP7_75t_R ALU___U645 ( .A(ALU__n773), .Y(ALU__n574) );
  BUFx12f_ASAP7_75t_R ALU___U646 ( .A(ALU__n702), .Y(ALU__n575) );
  BUFx12f_ASAP7_75t_R ALU___U647 ( .A(ALU__n542), .Y(ALU__n576) );
  INVx4_ASAP7_75t_R ALU___U648 ( .A(ALU__n1416), .Y(ALU__n1301) );
  BUFx3_ASAP7_75t_R ALU___U649 ( .A(ALU__n578), .Y(ALU__n577) );
  BUFx2_ASAP7_75t_R ALU___U650 ( .A(ALU__n294), .Y(ALU__n578) );
  AO22x2_ASAP7_75t_R ALU___U651 ( .A1(ALU__N155), .A2(ALU__n1563), .B1(ALU__N264), .B2(ALU__n27), .Y(
        n294) );
  BUFx4f_ASAP7_75t_R ALU___U652 ( .A(ALU__n577), .Y(ALU__n664) );
  BUFx2_ASAP7_75t_R ALU___U653 ( .A(ALU__n212), .Y(ALU__n579) );
  INVx6_ASAP7_75t_R ALU___U654 ( .A(ALU__n1300), .Y(ALU__n1394) );
  BUFx2_ASAP7_75t_R ALU___U655 ( .A(ALU__n248), .Y(ALU__n580) );
  INVx6_ASAP7_75t_R ALU___U656 ( .A(ALU__n628), .Y(ALU__n1014) );
  BUFx2_ASAP7_75t_R ALU___U657 ( .A(ALU__n290), .Y(ALU__n581) );
  BUFx2_ASAP7_75t_R ALU___U658 ( .A(ALU__n328), .Y(ALU__n582) );
  INVx5_ASAP7_75t_R ALU___U659 ( .A(ALU__n608), .Y(ALU__n1361) );
  BUFx3_ASAP7_75t_R ALU___U660 ( .A(ALU__n584), .Y(ALU__n583) );
  BUFx2_ASAP7_75t_R ALU___U661 ( .A(ALU__n1676), .Y(ALU__n584) );
  BUFx2_ASAP7_75t_R ALU___U662 ( .A(ALU__n891), .Y(ALU__n585) );
  AO221x1_ASAP7_75t_R ALU___U663 ( .A1(n1010), .A2(ALU__n1744), .B1(
        n1215), .B2(ALU__n938), .C(ALU__n890), .Y(ALU__n1676) );
  BUFx3_ASAP7_75t_R ALU___U664 ( .A(ALU__n587), .Y(ALU__n586) );
  BUFx2_ASAP7_75t_R ALU___U665 ( .A(ALU__n173), .Y(ALU__n587) );
  BUFx3_ASAP7_75t_R ALU___U666 ( .A(ALU__n589), .Y(ALU__n588) );
  BUFx2_ASAP7_75t_R ALU___U667 ( .A(ALU__n171), .Y(ALU__n589) );
  BUFx3_ASAP7_75t_R ALU___U668 ( .A(ALU__n591), .Y(ALU__n590) );
  BUFx2_ASAP7_75t_R ALU___U669 ( .A(ALU__n221), .Y(ALU__n591) );
  BUFx3_ASAP7_75t_R ALU___U670 ( .A(ALU__n593), .Y(ALU__n592) );
  BUFx2_ASAP7_75t_R ALU___U671 ( .A(ALU__n219), .Y(ALU__n593) );
  BUFx3_ASAP7_75t_R ALU___U672 ( .A(ALU__n595), .Y(ALU__n594) );
  BUFx2_ASAP7_75t_R ALU___U673 ( .A(ALU__n257), .Y(ALU__n595) );
  BUFx3_ASAP7_75t_R ALU___U674 ( .A(ALU__n597), .Y(ALU__n596) );
  BUFx2_ASAP7_75t_R ALU___U675 ( .A(ALU__n255), .Y(ALU__n597) );
  AO22x2_ASAP7_75t_R ALU___U676 ( .A1(ALU__N302), .A2(ALU__n1516), .B1(ALU__N334), .B2(ALU__n1504), .Y(
        n256) );
  BUFx3_ASAP7_75t_R ALU___U677 ( .A(ALU__n599), .Y(ALU__n598) );
  BUFx2_ASAP7_75t_R ALU___U678 ( .A(ALU__n317), .Y(ALU__n599) );
  BUFx3_ASAP7_75t_R ALU___U679 ( .A(ALU__n601), .Y(ALU__n600) );
  BUFx2_ASAP7_75t_R ALU___U680 ( .A(ALU__n315), .Y(ALU__n601) );
  INVx4_ASAP7_75t_R ALU___U681 ( .A(ALU__n1406), .Y(ALU__n602) );
  CKINVDCx11_ASAP7_75t_R ALU___U682 ( .A(ALU__n1734), .Y(ALU__n1406) );
  BUFx4f_ASAP7_75t_R ALU___U683 ( .A(ALU__n604), .Y(ALU__n603) );
  BUFx3_ASAP7_75t_R ALU___U684 ( .A(ALU__n567), .Y(ALU__n604) );
  AO22x2_ASAP7_75t_R ALU___U685 ( .A1(ALU__N173), .A2(ALU__n1564), .B1(ALU__N282), .B2(ALU__n1535), .Y(
        n186) );
  INVx2_ASAP7_75t_R ALU___U686 ( .A(ALU__n138), .Y(ALU__n605) );
  BUFx2_ASAP7_75t_R ALU___U687 ( .A(ALU__n327), .Y(ALU__n606) );
  BUFx2_ASAP7_75t_R ALU___U688 ( .A(ALU__n1647), .Y(ALU__n607) );
  BUFx12f_ASAP7_75t_R ALU___U689 ( .A(ALU__n1760), .Y(ALU__n608) );
  BUFx12f_ASAP7_75t_R ALU___U690 ( .A(ALU__n1758), .Y(ALU__n609) );
  BUFx12f_ASAP7_75t_R ALU___U691 ( .A(ALU__n630), .Y(ALU__n610) );
  INVx4_ASAP7_75t_R ALU___U692 ( .A(ALU__n780), .Y(ALU__n1747) );
  BUFx12f_ASAP7_75t_R ALU___U693 ( .A(ALU__n612), .Y(ALU__n611) );
  BUFx12f_ASAP7_75t_R ALU___U694 ( .A(ALU__n1495), .Y(ALU__n612) );
  CKINVDCx5p33_ASAP7_75t_R ALU___U695 ( .A(ALU__n611), .Y(ALU__n1473) );
  BUFx12f_ASAP7_75t_R ALU___U696 ( .A(ALU__n1129), .Y(ALU__n1495) );
  BUFx2_ASAP7_75t_R ALU___U697 ( .A(ALU__n140), .Y(ALU__n613) );
  BUFx16f_ASAP7_75t_R ALU___U698 ( .A(ALU__n1453), .Y(ALU__n614) );
  BUFx12f_ASAP7_75t_R ALU___U699 ( .A(ALU__n1019), .Y(ALU__n1453) );
  BUFx6f_ASAP7_75t_R ALU___U700 ( .A(ALU__n1020), .Y(ALU__n1019) );
  BUFx4f_ASAP7_75t_R ALU___U701 ( .A(ALU__n490), .Y(ALU__n1020) );
  BUFx3_ASAP7_75t_R ALU___U702 ( .A(ALU__n616), .Y(ALU__n615) );
  BUFx2_ASAP7_75t_R ALU___U703 ( .A(ALU__n239), .Y(ALU__n616) );
  BUFx3_ASAP7_75t_R ALU___U704 ( .A(ALU__n618), .Y(ALU__n617) );
  BUFx2_ASAP7_75t_R ALU___U705 ( .A(ALU__n237), .Y(ALU__n618) );
  BUFx2_ASAP7_75t_R ALU___U706 ( .A(ALU__n1673), .Y(ALU__n619) );
  BUFx2_ASAP7_75t_R ALU___U707 ( .A(ALU__n1671), .Y(ALU__n620) );
  BUFx3_ASAP7_75t_R ALU___U708 ( .A(ALU__n622), .Y(ALU__n621) );
  BUFx2_ASAP7_75t_R ALU___U709 ( .A(ALU__n1672), .Y(ALU__n622) );
  AO221x1_ASAP7_75t_R ALU___U710 ( .A1(n1100), .A2(ALU__n1066), .B1(ALU__n934), 
        .B2(ALU__n1687), .C(ALU__n620), .Y(ALU__n1672) );
  BUFx12f_ASAP7_75t_R ALU___U711 ( .A(ALU__n625), .Y(ALU__n623) );
  BUFx12f_ASAP7_75t_R ALU___U712 ( .A(ALU__n626), .Y(ALU__n624) );
  BUFx12f_ASAP7_75t_R ALU___U713 ( .A(ALU__n38), .Y(ALU__n625) );
  BUFx12f_ASAP7_75t_R ALU___U714 ( .A(ALU__n37), .Y(ALU__n626) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U715 ( .A(ALU__n624), .Y(ALU__n1600) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U716 ( .A(ALU__n623), .Y(ALU__n1601) );
  BUFx12f_ASAP7_75t_R ALU___U717 ( .A(ALU__n16), .Y(ALU__n776) );
  INVx2_ASAP7_75t_R ALU___U718 ( .A(ALU__n1548), .Y(ALU__n1529) );
  INVx2_ASAP7_75t_R ALU___U719 ( .A(ALU__n1582), .Y(ALU__n1557) );
  INVx4_ASAP7_75t_R ALU___U720 ( .A(n1056), .Y(ALU__n1689) );
  BUFx2_ASAP7_75t_R ALU___U721 ( .A(ALU__n246), .Y(ALU__n694) );
  INVx1_ASAP7_75t_R ALU___U722 ( .A(ALU__n694), .Y(ALU__n627) );
  BUFx12f_ASAP7_75t_R ALU___U723 ( .A(ALU__n1755), .Y(ALU__n628) );
  BUFx12f_ASAP7_75t_R ALU___U724 ( .A(ALU__n657), .Y(ALU__n629) );
  BUFx12f_ASAP7_75t_R ALU___U725 ( .A(ALU__n730), .Y(ALU__n630) );
  BUFx12f_ASAP7_75t_R ALU___U726 ( .A(ALU__n633), .Y(ALU__n631) );
  BUFx12f_ASAP7_75t_R ALU___U727 ( .A(ALU__n634), .Y(ALU__n632) );
  BUFx12f_ASAP7_75t_R ALU___U728 ( .A(ALU__n1273), .Y(ALU__n633) );
  BUFx12f_ASAP7_75t_R ALU___U729 ( .A(ALU__n1273), .Y(ALU__n634) );
  BUFx3_ASAP7_75t_R ALU___U730 ( .A(ALU__n636), .Y(ALU__n635) );
  BUFx2_ASAP7_75t_R ALU___U731 ( .A(ALU__n240), .Y(ALU__n636) );
  BUFx4f_ASAP7_75t_R ALU___U732 ( .A(ALU__n635), .Y(ALU__n689) );
  BUFx4f_ASAP7_75t_R ALU___U733 ( .A(ALU__n638), .Y(ALU__n637) );
  INVx2_ASAP7_75t_R ALU___U734 ( .A(ALU__n637), .Y(ALU__n1217) );
  BUFx4f_ASAP7_75t_R ALU___U735 ( .A(ALU__n1162), .Y(ALU__n639) );
  BUFx2_ASAP7_75t_R ALU___U736 ( .A(ALU__n139), .Y(ALU__n640) );
  INVx5_ASAP7_75t_R ALU___U737 ( .A(ALU__n1417), .Y(ALU__n1198) );
  BUFx4f_ASAP7_75t_R ALU___U738 ( .A(ALU__n642), .Y(ALU__n641) );
  BUFx3_ASAP7_75t_R ALU___U739 ( .A(ALU__n443), .Y(ALU__n642) );
  AO22x1_ASAP7_75t_R ALU___U740 ( .A1(ALU__N153), .A2(ALU__n1557), .B1(ALU__N262), .B2(ALU__n1526), .Y(
        n306) );
  BUFx2_ASAP7_75t_R ALU___U741 ( .A(ALU__n253), .Y(ALU__n643) );
  INVx5_ASAP7_75t_R ALU___U742 ( .A(ALU__n682), .Y(ALU__n982) );
  BUFx2_ASAP7_75t_R ALU___U743 ( .A(ALU__n325), .Y(ALU__n644) );
  BUFx12f_ASAP7_75t_R ALU___U744 ( .A(n422), .Y(ALU__n645) );
  BUFx12f_ASAP7_75t_R ALU___U745 ( .A(ALU__n602), .Y(ALU__n646) );
  BUFx16f_ASAP7_75t_R ALU___U746 ( .A(ALU__n645), .Y(ALU__n1734) );
  BUFx12f_ASAP7_75t_R ALU___U747 ( .A(ALU__n351), .Y(ALU__n648) );
  BUFx12f_ASAP7_75t_R ALU___U748 ( .A(ALU__n1521), .Y(ALU__n649) );
  BUFx12f_ASAP7_75t_R ALU___U749 ( .A(ALU__n743), .Y(ALU__n1521) );
  BUFx12f_ASAP7_75t_R ALU___U750 ( .A(ALU__n1364), .Y(ALU__n652) );
  BUFx12f_ASAP7_75t_R ALU___U751 ( .A(ALU__n1294), .Y(ALU__n1364) );
  AO22x2_ASAP7_75t_R ALU___U752 ( .A1(ALU__N179), .A2(ALU__n1567), .B1(ALU__N288), .B2(ALU__n1537), .Y(
        n150) );
  INVx2_ASAP7_75t_R ALU___U753 ( .A(ALU__n565), .Y(ALU__n653) );
  AO22x2_ASAP7_75t_R ALU___U754 ( .A1(ALU__N167), .A2(ALU__n1562), .B1(ALU__N276), .B2(ALU__n1532), .Y(
        n222) );
  INVx2_ASAP7_75t_R ALU___U755 ( .A(ALU__n403), .Y(ALU__n654) );
  BUFx2_ASAP7_75t_R ALU___U756 ( .A(ALU__n122), .Y(ALU__n655) );
  BUFx2_ASAP7_75t_R ALU___U757 ( .A(ALU__n1084), .Y(ALU__n656) );
  BUFx12f_ASAP7_75t_R ALU___U758 ( .A(ALU__n793), .Y(ALU__n657) );
  BUFx12f_ASAP7_75t_R ALU___U759 ( .A(ALU__n970), .Y(ALU__n658) );
  BUFx12f_ASAP7_75t_R ALU___U760 ( .A(ALU__n1448), .Y(ALU__n659) );
  CKINVDCx5p33_ASAP7_75t_R ALU___U761 ( .A(ALU__n1494), .Y(ALU__n1474) );
  BUFx12f_ASAP7_75t_R ALU___U762 ( .A(ALU__n1129), .Y(ALU__n1494) );
  AND2x4_ASAP7_75t_R ALU___U763 ( .A(ALU__N165), .B(ALU__n1561), .Y(ALU__n720) );
  INVx1_ASAP7_75t_R ALU___U764 ( .A(ALU__n720), .Y(ALU__n660) );
  AND2x4_ASAP7_75t_R ALU___U765 ( .A(ALU__N274), .B(ALU__n1531), .Y(ALU__n719) );
  INVx1_ASAP7_75t_R ALU___U766 ( .A(ALU__n719), .Y(ALU__n661) );
  AND2x2_ASAP7_75t_R ALU___U767 ( .A(ALU__n661), .B(ALU__n660), .Y(ALU__n234) );
  BUFx4f_ASAP7_75t_R ALU___U768 ( .A(ALU__n664), .Y(ALU__n663) );
  INVx2_ASAP7_75t_R ALU___U769 ( .A(ALU__n663), .Y(ALU__n1293) );
  BUFx12f_ASAP7_75t_R ALU___U770 ( .A(n637), .Y(ALU__n665) );
  BUFx16f_ASAP7_75t_R ALU___U771 ( .A(n637), .Y(ALU__n666) );
  BUFx16f_ASAP7_75t_R ALU___U772 ( .A(n637), .Y(ALU__n667) );
  BUFx4f_ASAP7_75t_R ALU___U773 ( .A(ALU__n669), .Y(ALU__n668) );
  BUFx3_ASAP7_75t_R ALU___U774 ( .A(ALU__n493), .Y(ALU__n669) );
  BUFx3_ASAP7_75t_R ALU___U775 ( .A(ALU__n671), .Y(ALU__n670) );
  BUFx2_ASAP7_75t_R ALU___U776 ( .A(ALU__n1658), .Y(ALU__n671) );
  BUFx2_ASAP7_75t_R ALU___U777 ( .A(ALU__n1657), .Y(ALU__n672) );
  BUFx3_ASAP7_75t_R ALU___U778 ( .A(ALU__n674), .Y(ALU__n673) );
  BUFx2_ASAP7_75t_R ALU___U779 ( .A(ALU__n1656), .Y(ALU__n674) );
  AO221x1_ASAP7_75t_R ALU___U780 ( .A1(n1109), .A2(ALU__n1345), .B1(
        n1152), .B2(ALU__n1297), .C(ALU__n672), .Y(ALU__n1658) );
  AO221x1_ASAP7_75t_R ALU___U781 ( .A1(n1029), .A2(ALU__n903), .B1(
        n1229), .B2(ALU__n1005), .C(ALU__n405), .Y(ALU__n1656) );
  BUFx10_ASAP7_75t_R ALU___U782 ( .A(ALU__n1299), .Y(ALU__n743) );
  BUFx16f_ASAP7_75t_R ALU___U783 ( .A(ALU__n1626), .Y(ALU__n676) );
  BUFx12f_ASAP7_75t_R ALU___U784 ( .A(ALU__n1294), .Y(ALU__n1626) );
  BUFx12f_ASAP7_75t_R ALU___U785 ( .A(ALU__n679), .Y(ALU__n677) );
  BUFx12f_ASAP7_75t_R ALU___U786 ( .A(ALU__n680), .Y(ALU__n678) );
  BUFx12f_ASAP7_75t_R ALU___U787 ( .A(ALU__n32), .Y(ALU__n679) );
  BUFx12f_ASAP7_75t_R ALU___U788 ( .A(ALU__n33), .Y(ALU__n680) );
  BUFx12f_ASAP7_75t_R ALU___U789 ( .A(ALU__n1425), .Y(ALU__n1614) );
  INVx2_ASAP7_75t_R ALU___U790 ( .A(ALU__n101), .Y(ALU__n681) );
  BUFx12f_ASAP7_75t_R ALU___U791 ( .A(ALU__n1754), .Y(ALU__n682) );
  BUFx12f_ASAP7_75t_R ALU___U792 ( .A(ALU__n684), .Y(ALU__n683) );
  BUFx12f_ASAP7_75t_R ALU___U793 ( .A(ALU__n610), .Y(ALU__n684) );
  INVx3_ASAP7_75t_R ALU___U794 ( .A(n955), .Y(ALU__n1688) );
  BUFx12f_ASAP7_75t_R ALU___U795 ( .A(ALU__n759), .Y(ALU__n685) );
  BUFx12f_ASAP7_75t_R ALU___U796 ( .A(ALU__n1447), .Y(ALU__n686) );
  BUFx12f_ASAP7_75t_R ALU___U797 ( .A(ALU__n1770), .Y(ALU__n687) );
  BUFx4f_ASAP7_75t_R ALU___U798 ( .A(ALU__n689), .Y(ALU__n688) );
  INVx2_ASAP7_75t_R ALU___U799 ( .A(ALU__n688), .Y(ALU__n1131) );
  BUFx2_ASAP7_75t_R ALU___U800 ( .A(ALU__n121), .Y(ALU__n690) );
  OR2x2_ASAP7_75t_R ALU___U801 ( .A(n1010), .B(ALU__n1744), .Y(ALU__n1677) );
  INVx1_ASAP7_75t_R ALU___U802 ( .A(ALU__n506), .Y(ALU__n691) );
  AND2x4_ASAP7_75t_R ALU___U803 ( .A(ALU__N163), .B(ALU__n1560), .Y(ALU__n723) );
  INVx1_ASAP7_75t_R ALU___U804 ( .A(ALU__n723), .Y(ALU__n692) );
  AND2x4_ASAP7_75t_R ALU___U805 ( .A(ALU__N272), .B(ALU__n1530), .Y(ALU__n722) );
  INVx1_ASAP7_75t_R ALU___U806 ( .A(ALU__n722), .Y(ALU__n693) );
  AND2x2_ASAP7_75t_R ALU___U807 ( .A(ALU__n693), .B(ALU__n692), .Y(ALU__n246) );
  BUFx12f_ASAP7_75t_R ALU___U808 ( .A(ALU__n696), .Y(ALU__n695) );
  BUFx12f_ASAP7_75t_R ALU___U809 ( .A(ALU__n1501), .Y(ALU__n696) );
  BUFx4f_ASAP7_75t_R ALU___U810 ( .A(ALU__n699), .Y(ALU__n698) );
  BUFx3_ASAP7_75t_R ALU___U811 ( .A(ALU__n340), .Y(ALU__n699) );
  INVx6_ASAP7_75t_R ALU___U812 ( .A(ALU__n695), .Y(ALU__n1396) );
  CKINVDCx5p33_ASAP7_75t_R ALU___U813 ( .A(ALU__n1517), .Y(ALU__n700) );
  BUFx16f_ASAP7_75t_R ALU___U814 ( .A(ALU__n648), .Y(ALU__n701) );
  BUFx12f_ASAP7_75t_R ALU___U815 ( .A(n553), .Y(ALU__n702) );
  BUFx10_ASAP7_75t_R ALU___U816 ( .A(ALU__n129), .Y(ALU__n1627) );
  CKINVDCx10_ASAP7_75t_R ALU___U817 ( .A(ALU__n112), .Y(ALU__n1620) );
  CKINVDCx10_ASAP7_75t_R ALU___U818 ( .A(ALU__n91), .Y(ALU__n1623) );
  BUFx12f_ASAP7_75t_R ALU___U819 ( .A(ALU__n26), .Y(ALU__n705) );
  BUFx12f_ASAP7_75t_R ALU___U820 ( .A(ALU__n105), .Y(ALU__n1612) );
  INVx6_ASAP7_75t_R ALU___U821 ( .A(ALU__n856), .Y(ALU__n1592) );
  INVx6_ASAP7_75t_R ALU___U822 ( .A(ALU__n398), .Y(ALU__n1591) );
  AO22x2_ASAP7_75t_R ALU___U823 ( .A1(ALU__N154), .A2(ALU__n1568), .B1(ALU__N263), .B2(ALU__n1527), .Y(
        n300) );
  INVx2_ASAP7_75t_R ALU___U824 ( .A(ALU__n547), .Y(ALU__n706) );
  INVx2_ASAP7_75t_R ALU___U825 ( .A(ALU__n346), .Y(ALU__n707) );
  BUFx12f_ASAP7_75t_R ALU___U826 ( .A(ALU__n935), .Y(ALU__n1768) );
  BUFx12f_ASAP7_75t_R ALU___U827 ( .A(ALU__n1752), .Y(ALU__n708) );
  INVx3_ASAP7_75t_R ALU___U828 ( .A(ALU__n1641), .Y(ALU__n1633) );
  BUFx6f_ASAP7_75t_R ALU___U829 ( .A(ALU__n860), .Y(ALU__n1641) );
  BUFx12f_ASAP7_75t_R ALU___U830 ( .A(ALU__n756), .Y(ALU__n709) );
  BUFx12f_ASAP7_75t_R ALU___U831 ( .A(ALU__n712), .Y(ALU__n710) );
  BUFx12f_ASAP7_75t_R ALU___U832 ( .A(ALU__n713), .Y(ALU__n711) );
  BUFx12f_ASAP7_75t_R ALU___U833 ( .A(ALU__n1272), .Y(ALU__n712) );
  BUFx12f_ASAP7_75t_R ALU___U834 ( .A(ALU__n712), .Y(ALU__n713) );
  BUFx12f_ASAP7_75t_R ALU___U835 ( .A(ALU__n785), .Y(ALU__n714) );
  BUFx12f_ASAP7_75t_R ALU___U836 ( .A(ALU__n1287), .Y(ALU__n715) );
  BUFx2_ASAP7_75t_R ALU___U837 ( .A(ALU__N224), .Y(ALU__n716) );
  BUFx4f_ASAP7_75t_R ALU___U838 ( .A(ALU__n1051), .Y(ALU__n717) );
  AO21x1_ASAP7_75t_R ALU___U839 ( .A1(ALU__n717), .A2(n888), .B(ALU__n1048), .Y(
        N224) );
  BUFx2_ASAP7_75t_R ALU___U840 ( .A(ALU__n569), .Y(ALU__n718) );
  INVx3_ASAP7_75t_R ALU___U841 ( .A(ALU__n13), .Y(ALU__n1561) );
  INVx4_ASAP7_75t_R ALU___U842 ( .A(ALU__n1545), .Y(ALU__n1531) );
  BUFx2_ASAP7_75t_R ALU___U843 ( .A(ALU__n627), .Y(ALU__n721) );
  INVx3_ASAP7_75t_R ALU___U844 ( .A(ALU__n1577), .Y(ALU__n1560) );
  INVx4_ASAP7_75t_R ALU___U845 ( .A(ALU__n1546), .Y(ALU__n1530) );
  BUFx12f_ASAP7_75t_R ALU___U846 ( .A(ALU__n1778), .Y(ALU__n724) );
  INVx2_ASAP7_75t_R ALU___U847 ( .A(ALU__N145), .Y(ALU__n1705) );
  BUFx12f_ASAP7_75t_R ALU___U848 ( .A(ALU__n726), .Y(ALU__n725) );
  BUFx12f_ASAP7_75t_R ALU___U849 ( .A(ALU__n1109), .Y(ALU__n726) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U850 ( .A(ALU__n725), .Y(ALU__n1483) );
  BUFx12f_ASAP7_75t_R ALU___U851 ( .A(ALU__n1493), .Y(ALU__n1109) );
  BUFx2_ASAP7_75t_R ALU___U852 ( .A(ALU__n120), .Y(ALU__n727) );
  BUFx4f_ASAP7_75t_R ALU___U853 ( .A(ALU__n729), .Y(ALU__n728) );
  INVx2_ASAP7_75t_R ALU___U854 ( .A(ALU__n728), .Y(ALU__n1316) );
  BUFx12f_ASAP7_75t_R ALU___U855 ( .A(n960), .Y(ALU__n730) );
  BUFx12f_ASAP7_75t_R ALU___U856 ( .A(n960), .Y(ALU__n731) );
  BUFx2_ASAP7_75t_R ALU___U857 ( .A(ALU__n1669), .Y(ALU__n732) );
  BUFx3_ASAP7_75t_R ALU___U858 ( .A(ALU__n734), .Y(ALU__n733) );
  BUFx2_ASAP7_75t_R ALU___U859 ( .A(ALU__n1670), .Y(ALU__n734) );
  BUFx3_ASAP7_75t_R ALU___U860 ( .A(ALU__n736), .Y(ALU__n735) );
  BUFx2_ASAP7_75t_R ALU___U861 ( .A(ALU__n1668), .Y(ALU__n736) );
  AO221x1_ASAP7_75t_R ALU___U862 ( .A1(n1064), .A2(ALU__n1688), .B1(
        n1178), .B2(ALU__n1689), .C(ALU__n732), .Y(ALU__n1670) );
  AO221x1_ASAP7_75t_R ALU___U863 ( .A1(n1024), .A2(ALU__n1106), .B1(
        n1225), .B2(ALU__n1741), .C(ALU__n425), .Y(ALU__n1668) );
  BUFx2_ASAP7_75t_R ALU___U864 ( .A(ALU__n1649), .Y(ALU__n737) );
  BUFx2_ASAP7_75t_R ALU___U865 ( .A(ALU__n1646), .Y(ALU__n738) );
  BUFx3_ASAP7_75t_R ALU___U866 ( .A(ALU__n740), .Y(ALU__n739) );
  BUFx2_ASAP7_75t_R ALU___U867 ( .A(ALU__n1648), .Y(ALU__n740) );
  AO221x1_ASAP7_75t_R ALU___U868 ( .A1(ALU__n1030), .A2(ALU__n1683), .B1(n1015), 
        .B2(ALU__n1053), .C(ALU__n738), .Y(ALU__n1648) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U869 ( .A(ALU__n1515), .Y(ALU__n741) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U870 ( .A(ALU__n1518), .Y(ALU__n742) );
  BUFx16f_ASAP7_75t_R ALU___U871 ( .A(ALU__n742), .Y(ALU__n1523) );
  BUFx12f_ASAP7_75t_R ALU___U872 ( .A(ALU__n1613), .Y(ALU__n744) );
  BUFx12f_ASAP7_75t_R ALU___U873 ( .A(ALU__n1425), .Y(ALU__n746) );
  CKINVDCx8_ASAP7_75t_R ALU___U874 ( .A(ALU__n1588), .Y(ALU__n1425) );
  INVx2_ASAP7_75t_R ALU___U875 ( .A(ALU__n383), .Y(ALU__n747) );
  BUFx12f_ASAP7_75t_R ALU___U876 ( .A(ALU__n1774), .Y(ALU__n1417) );
  BUFx6f_ASAP7_75t_R ALU___U877 ( .A(n1010), .Y(ALU__n1774) );
  BUFx12f_ASAP7_75t_R ALU___U878 ( .A(ALU__n1766), .Y(ALU__n748) );
  BUFx12f_ASAP7_75t_R ALU___U879 ( .A(ALU__n1780), .Y(ALU__n749) );
  BUFx16f_ASAP7_75t_R ALU___U880 ( .A(ALU__n1459), .Y(ALU__n750) );
  BUFx2_ASAP7_75t_R ALU___U881 ( .A(ALU__n1459), .Y(ALU__n751) );
  BUFx2_ASAP7_75t_R ALU___U882 ( .A(ALU__n1459), .Y(ALU__n752) );
  BUFx2_ASAP7_75t_R ALU___U883 ( .A(ALU__n1459), .Y(ALU__n753) );
  BUFx2_ASAP7_75t_R ALU___U884 ( .A(ALU__n1783), .Y(ALU__n754) );
  BUFx4f_ASAP7_75t_R ALU___U885 ( .A(ALU__n1240), .Y(EX_ALU_result[31]) );
  BUFx3_ASAP7_75t_R ALU___U886 ( .A(ALU__n754), .Y(ALU__n1240) );
  BUFx12f_ASAP7_75t_R ALU___U887 ( .A(ALU__n786), .Y(ALU__n755) );
  BUFx12f_ASAP7_75t_R ALU___U888 ( .A(ALU__n1034), .Y(ALU__n756) );
  BUFx16f_ASAP7_75t_R ALU___U889 ( .A(ALU__n832), .Y(ALU__n757) );
  BUFx6f_ASAP7_75t_R ALU___U890 ( .A(ALU__n832), .Y(ALU__n758) );
  BUFx12f_ASAP7_75t_R ALU___U891 ( .A(ALU__n1031), .Y(ALU__n759) );
  BUFx12f_ASAP7_75t_R ALU___U892 ( .A(ALU__n462), .Y(ALU__n760) );
  BUFx12f_ASAP7_75t_R ALU___U893 ( .A(ALU__n461), .Y(ALU__n761) );
  BUFx12f_ASAP7_75t_R ALU___U894 ( .A(ALU__n1202), .Y(ALU__n762) );
  BUFx12f_ASAP7_75t_R ALU___U895 ( .A(ALU__n764), .Y(ALU__n763) );
  BUFx12f_ASAP7_75t_R ALU___U896 ( .A(ALU__n1296), .Y(ALU__n764) );
  CKINVDCx5p33_ASAP7_75t_R ALU___U897 ( .A(ALU__n763), .Y(ALU__n1471) );
  BUFx12f_ASAP7_75t_R ALU___U898 ( .A(ALU__n68), .Y(ALU__n1296) );
  BUFx12f_ASAP7_75t_R ALU___U899 ( .A(ALU__n1512), .Y(ALU__n1506) );
  INVx6_ASAP7_75t_R ALU___U900 ( .A(ALU__n1511), .Y(ALU__n1502) );
  BUFx2_ASAP7_75t_R ALU___U901 ( .A(ALU__n1663), .Y(ALU__n765) );
  BUFx3_ASAP7_75t_R ALU___U902 ( .A(ALU__n767), .Y(ALU__n766) );
  BUFx2_ASAP7_75t_R ALU___U903 ( .A(ALU__n1662), .Y(ALU__n767) );
  BUFx3_ASAP7_75t_R ALU___U904 ( .A(ALU__n769), .Y(ALU__n768) );
  BUFx2_ASAP7_75t_R ALU___U905 ( .A(ALU__n1664), .Y(ALU__n769) );
  AO221x1_ASAP7_75t_R ALU___U906 ( .A1(n1073), .A2(ALU__n1695), .B1(
        n925), .B2(ALU__n1216), .C(ALU__n846), .Y(ALU__n1662) );
  AO221x1_ASAP7_75t_R ALU___U907 ( .A1(n1182), .A2(ALU__n1693), .B1(ALU__n966), 
        .B2(ALU__n1694), .C(ALU__n765), .Y(ALU__n1664) );
  INVx5_ASAP7_75t_R ALU___U908 ( .A(ALU__n1522), .Y(ALU__n1516) );
  BUFx12f_ASAP7_75t_R ALU___U909 ( .A(ALU__n741), .Y(ALU__n1522) );
  BUFx12f_ASAP7_75t_R ALU___U910 ( .A(ALU__n666), .Y(ALU__n770) );
  BUFx12f_ASAP7_75t_R ALU___U911 ( .A(ALU__n667), .Y(ALU__n771) );
  BUFx12f_ASAP7_75t_R ALU___U912 ( .A(ALU__n573), .Y(ALU__n772) );
  BUFx12f_ASAP7_75t_R ALU___U913 ( .A(ALU__n665), .Y(ALU__n773) );
  BUFx12f_ASAP7_75t_R ALU___U914 ( .A(ALU__n486), .Y(ALU__n899) );
  BUFx12f_ASAP7_75t_R ALU___U915 ( .A(ALU__n770), .Y(ALU__n902) );
  INVx4_ASAP7_75t_R ALU___U916 ( .A(n1091), .Y(ALU__n1775) );
  CKINVDCx10_ASAP7_75t_R ALU___U917 ( .A(ALU__n1532), .Y(ALU__n774) );
  BUFx12f_ASAP7_75t_R ALU___U918 ( .A(ALU__n1271), .Y(ALU__n1555) );
  BUFx12f_ASAP7_75t_R ALU___U919 ( .A(ALU__n775), .Y(ALU__n1583) );
  BUFx12f_ASAP7_75t_R ALU___U920 ( .A(ALU__n1608), .Y(ALU__n777) );
  BUFx12f_ASAP7_75t_R ALU___U921 ( .A(ALU__n77), .Y(ALU__ALU__n778) );
  BUFx12f_ASAP7_75t_R ALU___U922 ( .A(ALU__n576), .Y(ALU__n780) );
  BUFx12f_ASAP7_75t_R ALU___U923 ( .A(ALU__n543), .Y(ALU__n781) );
  BUFx12f_ASAP7_75t_R ALU___U924 ( .A(n553), .Y(ALU__n782) );
  BUFx12f_ASAP7_75t_R ALU___U925 ( .A(n553), .Y(ALU__n783) );
  INVx4_ASAP7_75t_R ALU___U926 ( .A(n790), .Y(ALU__n1694) );
  BUFx12f_ASAP7_75t_R ALU___U927 ( .A(ALU__n1737), .Y(ALU__n784) );
  BUFx12f_ASAP7_75t_R ALU___U928 ( .A(ALU__n967), .Y(ALU__n785) );
  BUFx12f_ASAP7_75t_R ALU___U929 ( .A(ALU__n935), .Y(ALU__n786) );
  BUFx2_ASAP7_75t_R ALU___U930 ( .A(ALU__n188), .Y(ALU__n787) );
  BUFx2_ASAP7_75t_R ALU___U931 ( .A(ALU__n260), .Y(ALU__n788) );
  BUFx2_ASAP7_75t_R ALU___U932 ( .A(ALU__n284), .Y(ALU__n789) );
  BUFx2_ASAP7_75t_R ALU___U933 ( .A(ALU__n302), .Y(ALU__n790) );
  BUFx2_ASAP7_75t_R ALU___U934 ( .A(ALU__n792), .Y(ALU__n791) );
  BUFx2_ASAP7_75t_R ALU___U935 ( .A(ALU__n124), .Y(ALU__n792) );
  BUFx12f_ASAP7_75t_R ALU___U936 ( .A(n777), .Y(ALU__n793) );
  BUFx12f_ASAP7_75t_R ALU___U937 ( .A(n777), .Y(ALU__n794) );
  BUFx2_ASAP7_75t_R ALU___U938 ( .A(ALU__n145), .Y(ALU__n795) );
  BUFx2_ASAP7_75t_R ALU___U939 ( .A(ALU__n313), .Y(ALU__n796) );
  BUFx3_ASAP7_75t_R ALU___U940 ( .A(ALU__n798), .Y(ALU__n797) );
  BUFx2_ASAP7_75t_R ALU___U941 ( .A(ALU__n233), .Y(ALU__n798) );
  BUFx3_ASAP7_75t_R ALU___U942 ( .A(ALU__n800), .Y(ALU__n799) );
  BUFx2_ASAP7_75t_R ALU___U943 ( .A(ALU__n231), .Y(ALU__n800) );
  BUFx3_ASAP7_75t_R ALU___U944 ( .A(ALU__n802), .Y(ALU__n801) );
  BUFx2_ASAP7_75t_R ALU___U945 ( .A(ALU__n287), .Y(ALU__n802) );
  BUFx3_ASAP7_75t_R ALU___U946 ( .A(ALU__n804), .Y(ALU__n803) );
  BUFx2_ASAP7_75t_R ALU___U947 ( .A(ALU__n285), .Y(ALU__n804) );
  BUFx2_ASAP7_75t_R ALU___U948 ( .A(ALU__n205), .Y(ALU__n805) );
  BUFx2_ASAP7_75t_R ALU___U949 ( .A(ALU__n277), .Y(ALU__n806) );
  CKINVDCx10_ASAP7_75t_R ALU___U950 ( .A(ALU__n55), .Y(ALU__n809) );
  BUFx2_ASAP7_75t_R ALU___U951 ( .A(ALU__N383), .Y(ALU__n810) );
  OA221x2_ASAP7_75t_R ALU___U952 ( .A1(ALU__n1705), .A2(ALU__n1622), .B1(ALU__n1362), .B2(ALU__n1599), 
        .C(ALU__n837), .Y(ALU__n161) );
  INVx1_ASAP7_75t_R ALU___U953 ( .A(ALU__n369), .Y(ALU__n811) );
  BUFx2_ASAP7_75t_R ALU___U954 ( .A(ALU__n160), .Y(ALU__n812) );
  OA22x2_ASAP7_75t_R ALU___U955 ( .A1(ALU__n917), .A2(ALU__n1685), .B1(ALU__n410), .B2(ALU__n530), .Y(
        n159) );
  INVx1_ASAP7_75t_R ALU___U956 ( .A(ALU__n371), .Y(ALU__n813) );
  INVx2_ASAP7_75t_R ALU___U957 ( .A(ALU__n1709), .Y(ALU__n1311) );
  BUFx2_ASAP7_75t_R ALU___U958 ( .A(ALU__n170), .Y(ALU__n814) );
  BUFx2_ASAP7_75t_R ALU___U959 ( .A(ALU__n176), .Y(ALU__n815) );
  BUFx2_ASAP7_75t_R ALU___U960 ( .A(ALU__n224), .Y(ALU__n816) );
  BUFx2_ASAP7_75t_R ALU___U961 ( .A(ALU__n314), .Y(ALU__n817) );
  BUFx2_ASAP7_75t_R ALU___U962 ( .A(ALU__n236), .Y(ALU__n818) );
  BUFx2_ASAP7_75t_R ALU___U963 ( .A(ALU__n125), .Y(ALU__n819) );
  BUFx4f_ASAP7_75t_R ALU___U964 ( .A(ALU__n821), .Y(ALU__n820) );
  INVx2_ASAP7_75t_R ALU___U965 ( .A(ALU__n820), .Y(ALU__n1334) );
  BUFx2_ASAP7_75t_R ALU___U966 ( .A(ALU__n217), .Y(ALU__n822) );
  BUFx3_ASAP7_75t_R ALU___U967 ( .A(ALU__n824), .Y(ALU__n823) );
  BUFx2_ASAP7_75t_R ALU___U968 ( .A(ALU__n149), .Y(ALU__n824) );
  BUFx3_ASAP7_75t_R ALU___U969 ( .A(ALU__n826), .Y(ALU__n825) );
  BUFx2_ASAP7_75t_R ALU___U970 ( .A(ALU__n147), .Y(ALU__n826) );
  AO22x2_ASAP7_75t_R ALU___U971 ( .A1(ALU__N320), .A2(ALU__n1519), .B1(ALU__N352), .B2(ALU__n1502), .Y(
        n148) );
  BUFx3_ASAP7_75t_R ALU___U972 ( .A(ALU__n828), .Y(ALU__n827) );
  BUFx2_ASAP7_75t_R ALU___U973 ( .A(ALU__n293), .Y(ALU__n828) );
  BUFx3_ASAP7_75t_R ALU___U974 ( .A(ALU__n830), .Y(ALU__n829) );
  BUFx2_ASAP7_75t_R ALU___U975 ( .A(ALU__n291), .Y(ALU__n830) );
  BUFx2_ASAP7_75t_R ALU___U976 ( .A(ALU__n319), .Y(ALU__n831) );
  BUFx12f_ASAP7_75t_R ALU___U977 ( .A(n779), .Y(ALU__n832) );
  BUFx2_ASAP7_75t_R ALU___U978 ( .A(ALU__N377), .Y(ALU__n833) );
  OA221x2_ASAP7_75t_R ALU___U979 ( .A1(ALU__n1312), .A2(ALU__n1620), .B1(ALU__n1335), .B2(ALU__n1598), 
        .C(ALU__n1003), .Y(ALU__n197) );
  INVx1_ASAP7_75t_R ALU___U980 ( .A(ALU__n411), .Y(ALU__n834) );
  OA22x2_ASAP7_75t_R ALU___U981 ( .A1(ALU__n519), .A2(ALU__n1741), .B1(n1075), .B2(
        n1195), .Y(ALU__n195) );
  INVx1_ASAP7_75t_R ALU___U982 ( .A(ALU__n413), .Y(ALU__n835) );
  BUFx2_ASAP7_75t_R ALU___U983 ( .A(ALU__n196), .Y(ALU__n836) );
  BUFx12f_ASAP7_75t_R ALU___U984 ( .A(ALU__n1772), .Y(ALU__n838) );
  BUFx12f_ASAP7_75t_R ALU___U985 ( .A(n1238), .Y(ALU__n935) );
  INVx6_ASAP7_75t_R ALU___U986 ( .A(ALU__n1505), .Y(ALU__n839) );
  BUFx2_ASAP7_75t_R ALU___U987 ( .A(ALU__n1786), .Y(ALU__n840) );
  BUFx2_ASAP7_75t_R ALU___U988 ( .A(ALU__n1792), .Y(ALU__n841) );
  BUFx2_ASAP7_75t_R ALU___U989 ( .A(ALU__n1798), .Y(ALU__n842) );
  BUFx12f_ASAP7_75t_R ALU___U990 ( .A(ALU__n1686), .Y(ALU__n843) );
  INVx2_ASAP7_75t_R ALU___U991 ( .A(ALU__n1712), .Y(ALU__n1292) );
  BUFx16f_ASAP7_75t_R ALU___U992 ( .A(ALU__n1107), .Y(ALU__n844) );
  BUFx12f_ASAP7_75t_R ALU___U993 ( .A(ALU__n1449), .Y(ALU__n1107) );
  BUFx12f_ASAP7_75t_R ALU___U994 ( .A(ALU__n1767), .Y(ALU__n845) );
  BUFx2_ASAP7_75t_R ALU___U995 ( .A(ALU__n1661), .Y(ALU__n846) );
  BUFx2_ASAP7_75t_R ALU___U996 ( .A(ALU__n1659), .Y(ALU__n847) );
  BUFx3_ASAP7_75t_R ALU___U997 ( .A(ALU__n849), .Y(ALU__n848) );
  BUFx2_ASAP7_75t_R ALU___U998 ( .A(ALU__n1660), .Y(ALU__n849) );
  AO221x1_ASAP7_75t_R ALU___U999 ( .A1(n969), .A2(ALU__n1697), .B1(
        n1020), .B2(ALU__n1738), .C(ALU__n847), .Y(ALU__n1660) );
  BUFx12f_ASAP7_75t_R ALU___U1000 ( .A(ALU__n850), .Y(ALU__n1492) );
  BUFx12f_ASAP7_75t_R ALU___U1001 ( .A(ALU__n1258), .Y(ALU__n1256) );
  BUFx3_ASAP7_75t_R ALU___U1002 ( .A(ALU__n852), .Y(EX_ALU_result[19]) );
  BUFx2_ASAP7_75t_R ALU___U1003 ( .A(ALU__n1795), .Y(ALU__n852) );
  INVx3_ASAP7_75t_R ALU___U1004 ( .A(ALU__n1524), .Y(ALU__n1514) );
  BUFx6f_ASAP7_75t_R ALU___U1005 ( .A(ALU__n741), .Y(ALU__n1524) );
  CKINVDCx12_ASAP7_75t_R ALU___U1006 ( .A(ALU__n1534), .Y(ALU__n853) );
  BUFx16f_ASAP7_75t_R ALU___U1007 ( .A(ALU__n853), .Y(ALU__n1546) );
  BUFx16f_ASAP7_75t_R ALU___U1008 ( .A(ALU__n1550), .Y(ALU__n1549) );
  BUFx12f_ASAP7_75t_R ALU___U1009 ( .A(ALU__n853), .Y(ALU__n1552) );
  CKINVDCx10_ASAP7_75t_R ALU___U1010 ( .A(ALU__n56), .Y(ALU__n855) );
  BUFx12f_ASAP7_75t_R ALU___U1011 ( .A(ALU__n1610), .Y(ALU__n856) );
  BUFx12f_ASAP7_75t_R ALU___U1012 ( .A(ALU__n1610), .Y(ALU__n858) );
  INVx4_ASAP7_75t_R ALU___U1013 ( .A(ALU__n1597), .Y(ALU__n859) );
  CKINVDCx10_ASAP7_75t_R ALU___U1014 ( .A(ALU__n65), .Y(ALU__n1597) );
  BUFx12f_ASAP7_75t_R ALU___U1015 ( .A(ALU__n862), .Y(ALU__n860) );
  BUFx12f_ASAP7_75t_R ALU___U1016 ( .A(ALU__n863), .Y(ALU__n861) );
  BUFx12f_ASAP7_75t_R ALU___U1017 ( .A(ALU__n1128), .Y(ALU__n862) );
  BUFx12f_ASAP7_75t_R ALU___U1018 ( .A(ALU__n1128), .Y(ALU__n863) );
  INVx2_ASAP7_75t_R ALU___U1019 ( .A(ALU__n1718), .Y(ALU__n1353) );
  INVx2_ASAP7_75t_R ALU___U1020 ( .A(ALU__n1702), .Y(ALU__n1252) );
  BUFx4f_ASAP7_75t_R ALU___U1021 ( .A(ALU__N148), .Y(ALU__n1702) );
  BUFx2_ASAP7_75t_R ALU___U1022 ( .A(ALU__n865), .Y(ALU__n864) );
  BUFx2_ASAP7_75t_R ALU___U1023 ( .A(ALU__n296), .Y(ALU__n865) );
  BUFx2_ASAP7_75t_R ALU___U1024 ( .A(ALU__n230), .Y(ALU__n866) );
  OR2x2_ASAP7_75t_R ALU___U1025 ( .A(ALU__n1411), .B(ALU__n1412), .Y(ALU__n122) );
  INVx1_ASAP7_75t_R ALU___U1026 ( .A(ALU__n655), .Y(ALU__n867) );
  BUFx2_ASAP7_75t_R ALU___U1027 ( .A(ALU__n1413), .Y(ALU__n868) );
  BUFx2_ASAP7_75t_R ALU___U1028 ( .A(ALU__n1414), .Y(ALU__n869) );
  INVx1_ASAP7_75t_R ALU___U1029 ( .A(ALU__n868), .Y(ALU__n1411) );
  INVx1_ASAP7_75t_R ALU___U1030 ( .A(ALU__n869), .Y(ALU__n1412) );
  BUFx6f_ASAP7_75t_R ALU___U1031 ( .A(n1105), .Y(ALU__n1035) );
  BUFx4f_ASAP7_75t_R ALU___U1032 ( .A(ALU__n871), .Y(ALU__n870) );
  BUFx3_ASAP7_75t_R ALU___U1033 ( .A(ALU__n71), .Y(ALU__n871) );
  BUFx2_ASAP7_75t_R ALU___U1034 ( .A(ALU__n187), .Y(ALU__n872) );
  BUFx2_ASAP7_75t_R ALU___U1035 ( .A(ALU__n223), .Y(ALU__n873) );
  BUFx2_ASAP7_75t_R ALU___U1036 ( .A(ALU__n259), .Y(ALU__n874) );
  BUFx3_ASAP7_75t_R ALU___U1037 ( .A(ALU__n876), .Y(ALU__n875) );
  BUFx2_ASAP7_75t_R ALU___U1038 ( .A(ALU__n245), .Y(ALU__n876) );
  BUFx3_ASAP7_75t_R ALU___U1039 ( .A(ALU__n878), .Y(ALU__n877) );
  BUFx2_ASAP7_75t_R ALU___U1040 ( .A(ALU__n243), .Y(ALU__n878) );
  BUFx3_ASAP7_75t_R ALU___U1041 ( .A(ALU__n880), .Y(ALU__n879) );
  BUFx2_ASAP7_75t_R ALU___U1042 ( .A(ALU__n269), .Y(ALU__n880) );
  BUFx3_ASAP7_75t_R ALU___U1043 ( .A(ALU__n882), .Y(ALU__n881) );
  BUFx2_ASAP7_75t_R ALU___U1044 ( .A(ALU__n267), .Y(ALU__n882) );
  BUFx3_ASAP7_75t_R ALU___U1045 ( .A(ALU__n884), .Y(ALU__n883) );
  BUFx2_ASAP7_75t_R ALU___U1046 ( .A(ALU__n311), .Y(ALU__n884) );
  BUFx3_ASAP7_75t_R ALU___U1047 ( .A(ALU__n886), .Y(ALU__n885) );
  BUFx2_ASAP7_75t_R ALU___U1048 ( .A(ALU__n309), .Y(ALU__n886) );
  BUFx2_ASAP7_75t_R ALU___U1049 ( .A(ALU__n136), .Y(ALU__n887) );
  BUFx2_ASAP7_75t_R ALU___U1050 ( .A(ALU__n289), .Y(ALU__n888) );
  INVx5_ASAP7_75t_R ALU___U1051 ( .A(ALU__n1009), .Y(ALU__n1363) );
  BUFx12f_ASAP7_75t_R ALU___U1052 ( .A(ALU__n111), .Y(ALU__n1748) );
  BUFx2_ASAP7_75t_R ALU___U1053 ( .A(ALU__n156), .Y(ALU__n889) );
  AO22x2_ASAP7_75t_R ALU___U1054 ( .A1(ALU__N178), .A2(ALU__n1567), .B1(ALU__N287), .B2(ALU__n1537), .Y(
        n156) );
  BUFx2_ASAP7_75t_R ALU___U1055 ( .A(ALU__n1675), .Y(ALU__n890) );
  INVx1_ASAP7_75t_R ALU___U1056 ( .A(ALU__n583), .Y(ALU__n891) );
  BUFx3_ASAP7_75t_R ALU___U1057 ( .A(ALU__n893), .Y(ALU__n892) );
  BUFx2_ASAP7_75t_R ALU___U1058 ( .A(ALU__n1674), .Y(ALU__n893) );
  AO221x1_ASAP7_75t_R ALU___U1059 ( .A1(n920), .A2(ALU__n1105), .B1(
        n1160), .B2(ALU__n1685), .C(ALU__n619), .Y(ALU__n1674) );
  BUFx2_ASAP7_75t_R ALU___U1060 ( .A(ALU__N375), .Y(ALU__n894) );
  OA221x2_ASAP7_75t_R ALU___U1061 ( .A1(ALU__n1333), .A2(ALU__n1621), .B1(ALU__n1394), .B2(ALU__n1599), 
        .C(ALU__n937), .Y(ALU__n209) );
  INVx1_ASAP7_75t_R ALU___U1062 ( .A(ALU__n555), .Y(ALU__n895) );
  BUFx2_ASAP7_75t_R ALU___U1063 ( .A(ALU__n208), .Y(ALU__n896) );
  OA22x2_ASAP7_75t_R ALU___U1064 ( .A1(ALU__n979), .A2(ALU__n1298), .B1(ALU__n794), .B2(ALU__n579), .Y(
        n207) );
  INVx1_ASAP7_75t_R ALU___U1065 ( .A(ALU__n557), .Y(ALU__n897) );
  INVx2_ASAP7_75t_R ALU___U1066 ( .A(ALU__n109), .Y(ALU__n898) );
  INVx3_ASAP7_75t_R ALU___U1067 ( .A(n619), .Y(ALU__n1680) );
  BUFx12f_ASAP7_75t_R ALU___U1068 ( .A(ALU__n772), .Y(ALU__n900) );
  BUFx12f_ASAP7_75t_R ALU___U1069 ( .A(ALU__n771), .Y(ALU__n901) );
  BUFx6f_ASAP7_75t_R ALU___U1070 ( .A(ALU_ctl[1]), .Y(ALU__n1735) );
  INVx3_ASAP7_75t_R ALU___U1071 ( .A(ALU__n1735), .Y(ALU__n988) );
  BUFx6f_ASAP7_75t_R ALU___U1072 ( .A(n1208), .Y(ALU__n1750) );
  INVx4_ASAP7_75t_R ALU___U1073 ( .A(ALU__n1750), .Y(ALU__n903) );
  BUFx12f_ASAP7_75t_R ALU___U1074 ( .A(n1105), .Y(ALU__n904) );
  BUFx6f_ASAP7_75t_R ALU___U1075 ( .A(ALU__n1033), .Y(ALU__n905) );
  BUFx12f_ASAP7_75t_R ALU___U1076 ( .A(n1096), .Y(ALU__n1030) );
  BUFx12f_ASAP7_75t_R ALU___U1077 ( .A(n1096), .Y(ALU__n1032) );
  INVx2_ASAP7_75t_R ALU___U1078 ( .A(ALU__n1726), .Y(ALU__n1254) );
  BUFx4f_ASAP7_75t_R ALU___U1079 ( .A(ALU__N124), .Y(ALU__n1726) );
  BUFx12f_ASAP7_75t_R ALU___U1080 ( .A(ALU__n908), .Y(ALU__n906) );
  BUFx12f_ASAP7_75t_R ALU___U1081 ( .A(ALU__n908), .Y(ALU__n907) );
  BUFx12f_ASAP7_75t_R ALU___U1082 ( .A(ALU__n987), .Y(ALU__n908) );
  BUFx4f_ASAP7_75t_R ALU___U1083 ( .A(ALU__n984), .Y(ALU__n909) );
  BUFx2_ASAP7_75t_R ALU___U1084 ( .A(ALU__n1429), .Y(ALU__n910) );
  AND5x1_ASAP7_75t_R ALU___U1085 ( .A(ALU__n1463), .B(ALU__n1490), .C(ALU__n1520), .D(ALU__n1539), .E(
        n1430), .Y(ALU__n1429) );
  BUFx2_ASAP7_75t_R ALU___U1086 ( .A(ALU__n690), .Y(ALU__n911) );
  BUFx4f_ASAP7_75t_R ALU___U1087 ( .A(ALU__n913), .Y(ALU__n912) );
  BUFx3_ASAP7_75t_R ALU___U1088 ( .A(ALU__n718), .Y(ALU__n913) );
  BUFx4f_ASAP7_75t_R ALU___U1089 ( .A(ALU__n915), .Y(ALU__n914) );
  BUFx3_ASAP7_75t_R ALU___U1090 ( .A(ALU__n342), .Y(ALU__n915) );
  BUFx2_ASAP7_75t_R ALU___U1091 ( .A(ALU__n151), .Y(ALU__n916) );
  BUFx2_ASAP7_75t_R ALU___U1092 ( .A(ALU__n163), .Y(ALU__n917) );
  BUFx2_ASAP7_75t_R ALU___U1093 ( .A(ALU__n247), .Y(ALU__n918) );
  BUFx2_ASAP7_75t_R ALU___U1094 ( .A(ALU__n265), .Y(ALU__n919) );
  BUFx2_ASAP7_75t_R ALU___U1095 ( .A(ALU__n295), .Y(ALU__n920) );
  BUFx3_ASAP7_75t_R ALU___U1096 ( .A(ALU__n922), .Y(ALU__n921) );
  BUFx2_ASAP7_75t_R ALU___U1097 ( .A(ALU__n251), .Y(ALU__n922) );
  BUFx3_ASAP7_75t_R ALU___U1098 ( .A(ALU__n924), .Y(ALU__n923) );
  BUFx2_ASAP7_75t_R ALU___U1099 ( .A(ALU__n249), .Y(ALU__n924) );
  BUFx2_ASAP7_75t_R ALU___U1100 ( .A(ALU__n169), .Y(ALU__n925) );
  INVx5_ASAP7_75t_R ALU___U1101 ( .A(ALU__n1236), .Y(ALU__n1419) );
  OR2x2_ASAP7_75t_R ALU___U1102 ( .A(ALU__n927), .B(ALU__n928), .Y(ALU__n137) );
  INVx1_ASAP7_75t_R ALU___U1103 ( .A(ALU__n469), .Y(ALU__n926) );
  OR2x2_ASAP7_75t_R ALU___U1104 ( .A(ALU__n1483), .B(ALU__n1775), .Y(ALU__n1407) );
  INVx1_ASAP7_75t_R ALU___U1105 ( .A(ALU__n471), .Y(ALU__n927) );
  OR2x2_ASAP7_75t_R ALU___U1106 ( .A(n1091), .B(ALU__n1454), .Y(ALU__n1408) );
  INVx1_ASAP7_75t_R ALU___U1107 ( .A(ALU__n472), .Y(ALU__n928) );
  AO22x2_ASAP7_75t_R ALU___U1108 ( .A1(ALU__N152), .A2(ALU__n1557), .B1(ALU__N261), .B2(ALU__n1526), .Y(
        n312) );
  INVx2_ASAP7_75t_R ALU___U1109 ( .A(ALU__n517), .Y(ALU__n929) );
  BUFx2_ASAP7_75t_R ALU___U1110 ( .A(ALU__N364), .Y(ALU__n930) );
  BUFx2_ASAP7_75t_R ALU___U1111 ( .A(ALU__n274), .Y(ALU__n931) );
  OA221x2_ASAP7_75t_R ALU___U1112 ( .A1(ALU__n1355), .A2(ALU__n1618), .B1(ALU__n1390), .B2(ALU__n1603), 
        .C(ALU__n1316), .Y(ALU__n275) );
  INVx1_ASAP7_75t_R ALU___U1113 ( .A(ALU__n438), .Y(ALU__n932) );
  OA22x2_ASAP7_75t_R ALU___U1114 ( .A1(ALU__n806), .A2(ALU__n1749), .B1(n619), .B2(
        n545), .Y(ALU__n273) );
  INVx1_ASAP7_75t_R ALU___U1115 ( .A(ALU__n440), .Y(ALU__n933) );
  BUFx12f_ASAP7_75t_R ALU___U1116 ( .A(n1238), .Y(ALU__n934) );
  BUFx12f_ASAP7_75t_R ALU___U1117 ( .A(n1238), .Y(ALU__n936) );
  BUFx6f_ASAP7_75t_R ALU___U1118 ( .A(n1123), .Y(ALU__n1684) );
  INVx4_ASAP7_75t_R ALU___U1119 ( .A(ALU__n1684), .Y(ALU__n938) );
  BUFx2_ASAP7_75t_R ALU___U1120 ( .A(ALU__n1805), .Y(ALU__n939) );
  BUFx12f_ASAP7_75t_R ALU___U1121 ( .A(ALU__n1036), .Y(ALU__n1761) );
  BUFx12f_ASAP7_75t_R ALU___U1122 ( .A(n1105), .Y(ALU__n1034) );
  BUFx12f_ASAP7_75t_R ALU___U1123 ( .A(ALU__n1757), .Y(ALU__n940) );
  INVx5_ASAP7_75t_R ALU___U1124 ( .A(ALU__n940), .Y(ALU__n1336) );
  BUFx4f_ASAP7_75t_R ALU___U1125 ( .A(ALU__n942), .Y(ALU__n941) );
  BUFx3_ASAP7_75t_R ALU___U1126 ( .A(ALU__n721), .Y(ALU__n942) );
  BUFx2_ASAP7_75t_R ALU___U1127 ( .A(ALU__n229), .Y(ALU__n943) );
  BUFx2_ASAP7_75t_R ALU___U1128 ( .A(ALU__n283), .Y(ALU__n944) );
  BUFx3_ASAP7_75t_R ALU___U1129 ( .A(ALU__n946), .Y(ALU__n945) );
  BUFx2_ASAP7_75t_R ALU___U1130 ( .A(ALU__n143), .Y(ALU__n946) );
  BUFx3_ASAP7_75t_R ALU___U1131 ( .A(ALU__n948), .Y(ALU__n947) );
  BUFx2_ASAP7_75t_R ALU___U1132 ( .A(ALU__n141), .Y(ALU__n948) );
  BUFx3_ASAP7_75t_R ALU___U1133 ( .A(ALU__n950), .Y(ALU__n949) );
  BUFx2_ASAP7_75t_R ALU___U1134 ( .A(ALU__n263), .Y(ALU__n950) );
  BUFx3_ASAP7_75t_R ALU___U1135 ( .A(ALU__n952), .Y(ALU__n951) );
  BUFx2_ASAP7_75t_R ALU___U1136 ( .A(ALU__n261), .Y(ALU__n952) );
  BUFx2_ASAP7_75t_R ALU___U1137 ( .A(ALU__n193), .Y(ALU__n953) );
  BUFx3_ASAP7_75t_R ALU___U1138 ( .A(ALU__n955), .Y(EX_ALU_result[12]) );
  BUFx2_ASAP7_75t_R ALU___U1139 ( .A(ALU__n1802), .Y(ALU__n955) );
  NOR2x1p5_ASAP7_75t_R ALU___U1140 ( .A(ALU_ctl[1]), .B(ALU__n1349), .Y(ALU__n1428) );
  BUFx4f_ASAP7_75t_R ALU___U1141 ( .A(ALU__n957), .Y(ALU__n956) );
  BUFx3_ASAP7_75t_R ALU___U1142 ( .A(ALU__n889), .Y(ALU__n957) );
  AO22x2_ASAP7_75t_R ALU___U1143 ( .A1(ALU__N161), .A2(ALU__n1566), .B1(ALU__N270), .B2(ALU__n1538), .Y(
        n258) );
  INVx2_ASAP7_75t_R ALU___U1144 ( .A(ALU__n914), .Y(ALU__n958) );
  AO22x2_ASAP7_75t_R ALU___U1145 ( .A1(ALU__N151), .A2(ALU__n1556), .B1(ALU__N260), .B2(ALU__n1525), .Y(
        n318) );
  INVx2_ASAP7_75t_R ALU___U1146 ( .A(ALU__n549), .Y(ALU__n959) );
  INVx2_ASAP7_75t_R ALU___U1147 ( .A(ALU__n641), .Y(ALU__n960) );
  BUFx2_ASAP7_75t_R ALU___U1148 ( .A(ALU__N362), .Y(ALU__n961) );
  BUFx2_ASAP7_75t_R ALU___U1149 ( .A(ALU__n286), .Y(ALU__n962) );
  OA221x2_ASAP7_75t_R ALU___U1150 ( .A1(ALU__n1254), .A2(ALU__n1623), .B1(ALU__n1363), .B2(ALU__n1602), 
        .C(ALU__n1132), .Y(ALU__n287) );
  INVx1_ASAP7_75t_R ALU___U1151 ( .A(ALU__n801), .Y(ALU__n963) );
  OA22x2_ASAP7_75t_R ALU___U1152 ( .A1(ALU__n888), .A2(ALU__n1194), .B1(ALU__n73), .B2(ALU__n581), .Y(
        n285) );
  INVx1_ASAP7_75t_R ALU___U1153 ( .A(ALU__n803), .Y(ALU__n964) );
  BUFx12f_ASAP7_75t_R ALU___U1154 ( .A(n1243), .Y(ALU__n965) );
  BUFx12f_ASAP7_75t_R ALU___U1155 ( .A(n1243), .Y(ALU__n966) );
  BUFx12f_ASAP7_75t_R ALU___U1156 ( .A(n1243), .Y(ALU__n967) );
  BUFx12f_ASAP7_75t_R ALU___U1157 ( .A(n1243), .Y(ALU__n968) );
  BUFx12f_ASAP7_75t_R ALU___U1158 ( .A(ALU__n757), .Y(ALU__n969) );
  BUFx12f_ASAP7_75t_R ALU___U1159 ( .A(n779), .Y(ALU__n970) );
  BUFx12f_ASAP7_75t_R ALU___U1160 ( .A(n779), .Y(ALU__n971) );
  BUFx2_ASAP7_75t_R ALU___U1161 ( .A(ALU__n727), .Y(ALU__n972) );
  BUFx12f_ASAP7_75t_R ALU___U1162 ( .A(n964), .Y(ALU__n1751) );
  BUFx2_ASAP7_75t_R ALU___U1163 ( .A(ALU__n175), .Y(ALU__n973) );
  BUFx2_ASAP7_75t_R ALU___U1164 ( .A(ALU__n235), .Y(ALU__n974) );
  BUFx3_ASAP7_75t_R ALU___U1165 ( .A(ALU__n976), .Y(ALU__n975) );
  BUFx2_ASAP7_75t_R ALU___U1166 ( .A(ALU__n179), .Y(ALU__n976) );
  BUFx3_ASAP7_75t_R ALU___U1167 ( .A(ALU__n978), .Y(ALU__n977) );
  BUFx2_ASAP7_75t_R ALU___U1168 ( .A(ALU__n177), .Y(ALU__n978) );
  INVx1_ASAP7_75t_R ALU___U1169 ( .A(n955), .Y(ALU__n1742) );
  BUFx2_ASAP7_75t_R ALU___U1170 ( .A(ALU__n211), .Y(ALU__n979) );
  BUFx2_ASAP7_75t_R ALU___U1171 ( .A(ALU__n271), .Y(ALU__n980) );
  INVx5_ASAP7_75t_R ALU___U1172 ( .A(ALU__n1238), .Y(ALU__n1389) );
  BUFx12f_ASAP7_75t_R ALU___U1173 ( .A(ALU__n62), .Y(ALU__n1699) );
  BUFx12f_ASAP7_75t_R ALU___U1174 ( .A(ALU__n51), .Y(ALU__n1681) );
  BUFx6f_ASAP7_75t_R ALU___U1175 ( .A(n1073), .Y(ALU__n1758) );
  BUFx6f_ASAP7_75t_R ALU___U1176 ( .A(n1109), .Y(ALU__n1754) );
  BUFx6f_ASAP7_75t_R ALU___U1177 ( .A(ALU__n909), .Y(ALU__n983) );
  BUFx3_ASAP7_75t_R ALU___U1178 ( .A(ALU__n910), .Y(ALU__n984) );
  BUFx12f_ASAP7_75t_R ALU___U1179 ( .A(ALU__n907), .Y(ALU__n985) );
  BUFx12f_ASAP7_75t_R ALU___U1180 ( .A(ALU__n906), .Y(ALU__n986) );
  BUFx12f_ASAP7_75t_R ALU___U1181 ( .A(ALU__n1645), .Y(ALU__n987) );
  BUFx12f_ASAP7_75t_R ALU___U1182 ( .A(ALU__n983), .Y(ALU__n1645) );
  AO22x2_ASAP7_75t_R ALU___U1183 ( .A1(ALU__N160), .A2(ALU__n1565), .B1(ALU__N269), .B2(ALU__n1533), .Y(
        n264) );
  INVx2_ASAP7_75t_R ALU___U1184 ( .A(ALU__n870), .Y(ALU__n989) );
  INVx2_ASAP7_75t_R ALU___U1185 ( .A(ALU__n956), .Y(ALU__n990) );
  BUFx2_ASAP7_75t_R ALU___U1186 ( .A(ALU__N386), .Y(ALU__n991) );
  OA221x2_ASAP7_75t_R ALU___U1187 ( .A1(ALU__n1252), .A2(ALU__n1623), .B1(ALU__n1198), .B2(ALU__n1603), 
        .C(ALU__n1063), .Y(ALU__n143) );
  INVx1_ASAP7_75t_R ALU___U1188 ( .A(ALU__n945), .Y(ALU__n992) );
  BUFx2_ASAP7_75t_R ALU___U1189 ( .A(ALU__n142), .Y(ALU__n993) );
  OA22x2_ASAP7_75t_R ALU___U1190 ( .A1(ALU__n795), .A2(ALU__n1744), .B1(ALU__n731), .B2(ALU__n442), .Y(
        n141) );
  INVx1_ASAP7_75t_R ALU___U1191 ( .A(ALU__n947), .Y(ALU__n994) );
  BUFx2_ASAP7_75t_R ALU___U1192 ( .A(ALU__N374), .Y(ALU__n995) );
  OA221x2_ASAP7_75t_R ALU___U1193 ( .A1(ALU__n1329), .A2(ALU__n1622), .B1(ALU__n1361), .B2(ALU__n1599), 
        .C(ALU__n747), .Y(ALU__n215) );
  INVx1_ASAP7_75t_R ALU___U1194 ( .A(ALU__n448), .Y(ALU__n996) );
  OA22x2_ASAP7_75t_R ALU___U1195 ( .A1(ALU__n822), .A2(ALU__n1693), .B1(n858), 
        .B2(ALU__n531), .Y(ALU__n213) );
  INVx1_ASAP7_75t_R ALU___U1196 ( .A(ALU__n450), .Y(ALU__n997) );
  BUFx2_ASAP7_75t_R ALU___U1197 ( .A(ALU__n214), .Y(ALU__n998) );
  BUFx2_ASAP7_75t_R ALU___U1198 ( .A(ALU__N358), .Y(ALU__n999) );
  BUFx2_ASAP7_75t_R ALU___U1199 ( .A(ALU__n310), .Y(ALU__n1000) );
  OA221x2_ASAP7_75t_R ALU___U1200 ( .A1(ALU__n1377), .A2(ALU__n1623), .B1(ALU__n1301), .B2(ALU__n1604), 
        .C(ALU__n929), .Y(ALU__n311) );
  INVx1_ASAP7_75t_R ALU___U1201 ( .A(ALU__n883), .Y(ALU__n1001) );
  OA22x2_ASAP7_75t_R ALU___U1202 ( .A1(ALU__n796), .A2(ALU__n484), .B1(ALU__n969), .B2(ALU__n817), .Y(
        n309) );
  INVx1_ASAP7_75t_R ALU___U1203 ( .A(ALU__n885), .Y(ALU__n1002) );
  BUFx2_ASAP7_75t_R ALU___U1204 ( .A(ALU__n1809), .Y(ALU__n1004) );
  BUFx4f_ASAP7_75t_R ALU___U1205 ( .A(ALU__n1207), .Y(EX_ALU_result[5]) );
  BUFx3_ASAP7_75t_R ALU___U1206 ( .A(ALU__n1004), .Y(ALU__n1207) );
  BUFx6f_ASAP7_75t_R ALU___U1207 ( .A(n1164), .Y(ALU__n1737) );
  INVx4_ASAP7_75t_R ALU___U1208 ( .A(ALU__n784), .Y(ALU__n1005) );
  BUFx2_ASAP7_75t_R ALU___U1209 ( .A(ALU__n1784), .Y(ALU__n1006) );
  BUFx2_ASAP7_75t_R ALU___U1210 ( .A(ALU__n1806), .Y(ALU__n1007) );
  INVx2_ASAP7_75t_R ALU___U1211 ( .A(ALU__n1721), .Y(ALU__n1317) );
  BUFx2_ASAP7_75t_R ALU___U1212 ( .A(ALU__n158), .Y(ALU__n1008) );
  BUFx12f_ASAP7_75t_R ALU___U1213 ( .A(ALU__n1779), .Y(ALU__n1009) );
  BUFx3_ASAP7_75t_R ALU___U1214 ( .A(ALU__n1011), .Y(ALU__n1010) );
  BUFx2_ASAP7_75t_R ALU___U1215 ( .A(ALU__n203), .Y(ALU__n1011) );
  BUFx3_ASAP7_75t_R ALU___U1216 ( .A(ALU__n1013), .Y(ALU__n1012) );
  BUFx2_ASAP7_75t_R ALU___U1217 ( .A(ALU__n201), .Y(ALU__n1013) );
  BUFx6f_ASAP7_75t_R ALU___U1218 ( .A(n1020), .Y(ALU__n1755) );
  BUFx12f_ASAP7_75t_R ALU___U1219 ( .A(ALU__n1339), .Y(ALU__n1015) );
  BUFx12f_ASAP7_75t_R ALU___U1220 ( .A(ALU__n42), .Y(ALU__n1339) );
  BUFx3_ASAP7_75t_R ALU___U1221 ( .A(ALU__n1017), .Y(EX_ALU_result[17]) );
  BUFx2_ASAP7_75t_R ALU___U1222 ( .A(ALU__n1797), .Y(ALU__n1017) );
  INVx3_ASAP7_75t_R ALU___U1223 ( .A(ALU__n1018), .Y(ALU__n1439) );
  OR3x1_ASAP7_75t_R ALU___U1224 ( .A(ALU_ctl[3]), .B(ALU__n646), .C(ALU_ctl[1]), 
        .Y(ALU__n140) );
  BUFx2_ASAP7_75t_R ALU___U1225 ( .A(ALU__n529), .Y(ALU__n324) );
  INVx2_ASAP7_75t_R ALU___U1226 ( .A(ALU__n527), .Y(ALU__n1021) );
  AND2x4_ASAP7_75t_R ALU___U1227 ( .A(ALU__N150), .B(ALU__n1556), .Y(ALU__n1423) );
  INVx1_ASAP7_75t_R ALU___U1228 ( .A(ALU__n1423), .Y(ALU__n1022) );
  AND2x4_ASAP7_75t_R ALU___U1229 ( .A(ALU__N259), .B(ALU__n1525), .Y(ALU__n1424) );
  INVx1_ASAP7_75t_R ALU___U1230 ( .A(ALU__n1424), .Y(ALU__n1023) );
  AND2x2_ASAP7_75t_R ALU___U1231 ( .A(ALU__n1022), .B(ALU__n1023), .Y(ALU__n1422) );
  INVx2_ASAP7_75t_R ALU___U1232 ( .A(ALU__n912), .Y(ALU__n1025) );
  BUFx2_ASAP7_75t_R ALU___U1233 ( .A(ALU__N385), .Y(ALU__n1026) );
  BUFx2_ASAP7_75t_R ALU___U1234 ( .A(ALU__n148), .Y(ALU__n1027) );
  OA221x2_ASAP7_75t_R ALU___U1235 ( .A1(ALU__n1310), .A2(ALU__n1623), .B1(ALU__n1358), .B2(ALU__n1602), 
        .C(ALU__n653), .Y(ALU__n149) );
  INVx1_ASAP7_75t_R ALU___U1236 ( .A(ALU__n823), .Y(ALU__n1028) );
  OA22x2_ASAP7_75t_R ALU___U1237 ( .A1(ALU__n916), .A2(ALU__n938), .B1(n1123), .B2(
        n365), .Y(ALU__n147) );
  INVx1_ASAP7_75t_R ALU___U1238 ( .A(ALU__n825), .Y(ALU__n1029) );
  BUFx12f_ASAP7_75t_R ALU___U1239 ( .A(n1096), .Y(ALU__n1031) );
  BUFx12f_ASAP7_75t_R ALU___U1240 ( .A(n1096), .Y(ALU__n1033) );
  BUFx12f_ASAP7_75t_R ALU___U1241 ( .A(n1105), .Y(ALU__n1036) );
  BUFx12f_ASAP7_75t_R ALU___U1242 ( .A(n1105), .Y(ALU__n1037) );
  INVx2_ASAP7_75t_R ALU___U1243 ( .A(ALU__n603), .Y(ALU__n1038) );
  BUFx12f_ASAP7_75t_R ALU___U1244 ( .A(ALU__n570), .Y(ALU__n1039) );
  BUFx16f_ASAP7_75t_R ALU___U1245 ( .A(ALU__n1461), .Y(ALU__n1040) );
  BUFx2_ASAP7_75t_R ALU___U1246 ( .A(ALU__n1461), .Y(ALU__n1041) );
  BUFx2_ASAP7_75t_R ALU___U1247 ( .A(ALU__n1461), .Y(ALU__n1042) );
  BUFx2_ASAP7_75t_R ALU___U1248 ( .A(ALU__n1461), .Y(ALU__n1043) );
  BUFx2_ASAP7_75t_R ALU___U1249 ( .A(ALU__n1791), .Y(ALU__n1044) );
  BUFx2_ASAP7_75t_R ALU___U1250 ( .A(ALU__n1808), .Y(ALU__n1045) );
  BUFx2_ASAP7_75t_R ALU___U1251 ( .A(ALU__n1812), .Y(ALU__n1046) );
  BUFx2_ASAP7_75t_R ALU___U1252 ( .A(ALU__n326), .Y(ALU__n1047) );
  BUFx2_ASAP7_75t_R ALU___U1253 ( .A(ALU__n1678), .Y(ALU__n1048) );
  BUFx4f_ASAP7_75t_R ALU___U1254 ( .A(ALU__n1050), .Y(ALU__n1049) );
  BUFx3_ASAP7_75t_R ALU___U1255 ( .A(ALU__n716), .Y(ALU__n1050) );
  BUFx4f_ASAP7_75t_R ALU___U1256 ( .A(n1091), .Y(ALU__n1679) );
  INVx2_ASAP7_75t_R ALU___U1257 ( .A(ALU__n1679), .Y(ALU__n1051) );
  BUFx12f_ASAP7_75t_R ALU___U1258 ( .A(ALU__n1765), .Y(ALU__n1052) );
  INVx5_ASAP7_75t_R ALU___U1259 ( .A(ALU__n1052), .Y(ALU__n1393) );
  BUFx4f_ASAP7_75t_R ALU___U1260 ( .A(ALU__n1054), .Y(ALU__n1053) );
  BUFx3_ASAP7_75t_R ALU___U1261 ( .A(ALU__n607), .Y(ALU__n1054) );
  INVx4_ASAP7_75t_R ALU___U1262 ( .A(n1152), .Y(ALU__n1753) );
  BUFx3_ASAP7_75t_R ALU___U1263 ( .A(ALU__n1057), .Y(EX_ALU_result[1]) );
  BUFx2_ASAP7_75t_R ALU___U1264 ( .A(ALU__n1813), .Y(ALU__n1057) );
  BUFx12f_ASAP7_75t_R ALU___U1265 ( .A(ALU__n1789), .Y(ALU__n1058) );
  BUFx4f_ASAP7_75t_R ALU___U1266 ( .A(ALU__N149), .Y(ALU__n1701) );
  INVx3_ASAP7_75t_R ALU___U1267 ( .A(ALU_ctl[3]), .Y(ALU__n1733) );
  NOR2x1p5_ASAP7_75t_R ALU___U1268 ( .A(ALU_ctl[3]), .B(ALU_ctl[1]), .Y(
        n1398) );
  BUFx2_ASAP7_75t_R ALU___U1269 ( .A(ALU__N370), .Y(ALU__n1059) );
  BUFx2_ASAP7_75t_R ALU___U1270 ( .A(ALU__n238), .Y(ALU__n1060) );
  OA221x2_ASAP7_75t_R ALU___U1271 ( .A1(ALU__n1353), .A2(ALU__n1620), .B1(ALU__n1337), .B2(ALU__n1600), 
        .C(ALU__n1131), .Y(ALU__n239) );
  INVx1_ASAP7_75t_R ALU___U1272 ( .A(ALU__n615), .Y(ALU__n1061) );
  OA22x2_ASAP7_75t_R ALU___U1273 ( .A1(ALU__n564), .A2(ALU__n1739), .B1(n794), 
        .B2(ALU__n515), .Y(ALU__n237) );
  INVx1_ASAP7_75t_R ALU___U1274 ( .A(ALU__n617), .Y(ALU__n1062) );
  INVx1_ASAP7_75t_R ALU___U1275 ( .A(n794), .Y(ALU__n1739) );
  AO22x1_ASAP7_75t_R ALU___U1276 ( .A1(ALU__N180), .A2(ALU__n1568), .B1(ALU__N289), .B2(ALU__n1538), .Y(
        n144) );
  BUFx2_ASAP7_75t_R ALU___U1277 ( .A(ALU__n1810), .Y(ALU__n1064) );
  BUFx4f_ASAP7_75t_R ALU___U1278 ( .A(ALU__n1279), .Y(EX_ALU_result[4]) );
  BUFx3_ASAP7_75t_R ALU___U1279 ( .A(ALU__n1064), .Y(ALU__n1279) );
  INVx2_ASAP7_75t_R ALU___U1280 ( .A(n858), .Y(ALU__n1065) );
  BUFx4f_ASAP7_75t_R ALU___U1281 ( .A(n978), .Y(ALU__n1686) );
  INVx4_ASAP7_75t_R ALU___U1282 ( .A(ALU__n843), .Y(ALU__n1066) );
  BUFx12f_ASAP7_75t_R ALU___U1283 ( .A(ALU__n1446), .Y(ALU__n1067) );
  BUFx12f_ASAP7_75t_R ALU___U1284 ( .A(ALU__n1451), .Y(ALU__n1446) );
  BUFx2_ASAP7_75t_R ALU___U1285 ( .A(ALU__n1785), .Y(ALU__n1068) );
  BUFx2_ASAP7_75t_R ALU___U1286 ( .A(ALU__n1793), .Y(ALU__n1069) );
  BUFx2_ASAP7_75t_R ALU___U1287 ( .A(ALU__n1799), .Y(ALU__n1070) );
  BUFx2_ASAP7_75t_R ALU___U1288 ( .A(ALU__n1807), .Y(ALU__n1071) );
  BUFx12f_ASAP7_75t_R ALU___U1289 ( .A(ALU__n1771), .Y(ALU__n1072) );
  BUFx12f_ASAP7_75t_R ALU___U1290 ( .A(ALU__n1763), .Y(ALU__n1073) );
  INVx5_ASAP7_75t_R ALU___U1291 ( .A(ALU__n1073), .Y(ALU__n1418) );
  BUFx3_ASAP7_75t_R ALU___U1292 ( .A(ALU__n1075), .Y(EX_ALU_result[11]) );
  BUFx2_ASAP7_75t_R ALU___U1293 ( .A(ALU__n1803), .Y(ALU__n1075) );
  BUFx12f_ASAP7_75t_R ALU___U1294 ( .A(ALU__n1078), .Y(ALU__n1077) );
  BUFx12f_ASAP7_75t_R ALU___U1295 ( .A(ALU__n1496), .Y(ALU__n1078) );
  INVx6_ASAP7_75t_R ALU___U1296 ( .A(ALU__n1077), .Y(ALU__n1472) );
  BUFx12f_ASAP7_75t_R ALU___U1297 ( .A(ALU__n69), .Y(ALU__n1496) );
  BUFx12f_ASAP7_75t_R ALU___U1298 ( .A(ALU__n1787), .Y(ALU__n1079) );
  INVx2_ASAP7_75t_R ALU___U1299 ( .A(ALU__n941), .Y(ALU__n1082) );
  BUFx3_ASAP7_75t_R ALU___U1300 ( .A(ALU__n656), .Y(ALU__n1083) );
  BUFx2_ASAP7_75t_R ALU___U1301 ( .A(ALU__N118), .Y(ALU__n1732) );
  INVx1_ASAP7_75t_R ALU___U1302 ( .A(ALU__n1732), .Y(ALU__n1084) );
  BUFx2_ASAP7_75t_R ALU___U1303 ( .A(ALU__N381), .Y(ALU__n1085) );
  BUFx2_ASAP7_75t_R ALU___U1304 ( .A(ALU__n172), .Y(ALU__n1086) );
  OA221x2_ASAP7_75t_R ALU___U1305 ( .A1(ALU__n1350), .A2(ALU__n1622), .B1(ALU__n1385), .B2(ALU__n1597), 
        .C(ALU__n568), .Y(ALU__n173) );
  INVx1_ASAP7_75t_R ALU___U1306 ( .A(ALU__n586), .Y(ALU__n1087) );
  OA22x2_ASAP7_75t_R ALU___U1307 ( .A1(ALU__n973), .A2(ALU__n1687), .B1(n851), 
        .B2(ALU__n815), .Y(ALU__n171) );
  INVx1_ASAP7_75t_R ALU___U1308 ( .A(ALU__n588), .Y(ALU__n1088) );
  BUFx2_ASAP7_75t_R ALU___U1309 ( .A(ALU__N373), .Y(ALU__n1089) );
  OA221x2_ASAP7_75t_R ALU___U1310 ( .A1(ALU__n1330), .A2(ALU__n1621), .B1(ALU__n1388), .B2(ALU__n1600), 
        .C(ALU__n654), .Y(ALU__n221) );
  INVx1_ASAP7_75t_R ALU___U1311 ( .A(ALU__n590), .Y(ALU__n1090) );
  OA22x2_ASAP7_75t_R ALU___U1312 ( .A1(ALU__n873), .A2(ALU__n1694), .B1(n790), 
        .B2(ALU__n816), .Y(ALU__n219) );
  INVx1_ASAP7_75t_R ALU___U1313 ( .A(ALU__n592), .Y(ALU__n1091) );
  BUFx2_ASAP7_75t_R ALU___U1314 ( .A(ALU__n220), .Y(ALU__n1092) );
  BUFx2_ASAP7_75t_R ALU___U1315 ( .A(ALU__N368), .Y(ALU__n1093) );
  BUFx2_ASAP7_75t_R ALU___U1316 ( .A(ALU__n250), .Y(ALU__n1094) );
  OA221x2_ASAP7_75t_R ALU___U1317 ( .A1(ALU__n1314), .A2(ALU__n1619), .B1(ALU__n982), .B2(ALU__n1602), 
        .C(ALU__n1409), .Y(ALU__n251) );
  INVx1_ASAP7_75t_R ALU___U1318 ( .A(ALU__n921), .Y(ALU__n1095) );
  OA22x2_ASAP7_75t_R ALU___U1319 ( .A1(ALU__n643), .A2(ALU__n1345), .B1(n352), 
        .B2(ALU__n516), .Y(ALU__n249) );
  INVx1_ASAP7_75t_R ALU___U1320 ( .A(ALU__n923), .Y(ALU__n1096) );
  BUFx2_ASAP7_75t_R ALU___U1321 ( .A(ALU__N357), .Y(ALU__n1097) );
  BUFx2_ASAP7_75t_R ALU___U1322 ( .A(ALU__n316), .Y(ALU__n1098) );
  OA221x2_ASAP7_75t_R ALU___U1323 ( .A1(ALU__n1253), .A2(ALU__n1618), .B1(ALU__n1415), .B2(ALU__n1604), 
        .C(ALU__n959), .Y(ALU__n317) );
  INVx1_ASAP7_75t_R ALU___U1324 ( .A(ALU__n598), .Y(ALU__n1099) );
  OA22x2_ASAP7_75t_R ALU___U1325 ( .A1(ALU__n831), .A2(ALU__n1289), .B1(n749), .B2(
        n1197), .Y(ALU__n315) );
  INVx1_ASAP7_75t_R ALU___U1326 ( .A(ALU__n600), .Y(ALU__n1100) );
  INVx1_ASAP7_75t_R ALU___U1327 ( .A(n779), .Y(ALU__n1743) );
  INVx3_ASAP7_75t_R ALU___U1328 ( .A(ALU__n758), .Y(ALU__n1683) );
  BUFx6f_ASAP7_75t_R ALU___U1329 ( .A(n1222), .Y(ALU__n1696) );
  BUFx16f_ASAP7_75t_R ALU___U1330 ( .A(ALU__n1462), .Y(ALU__n1101) );
  BUFx2_ASAP7_75t_R ALU___U1331 ( .A(ALU__n1462), .Y(ALU__n1102) );
  BUFx2_ASAP7_75t_R ALU___U1332 ( .A(ALU__n1462), .Y(ALU__n1103) );
  BUFx2_ASAP7_75t_R ALU___U1333 ( .A(ALU__n1462), .Y(ALU__n1104) );
  INVx4_ASAP7_75t_R ALU___U1334 ( .A(n1033), .Y(ALU__n1105) );
  INVx4_ASAP7_75t_R ALU___U1335 ( .A(n1162), .Y(ALU__n1106) );
  INVx2_ASAP7_75t_R ALU___U1336 ( .A(ALU__n1725), .Y(ALU__n1315) );
  INVx2_ASAP7_75t_R ALU___U1337 ( .A(ALU__n1729), .Y(ALU__n1354) );
  INVx2_ASAP7_75t_R ALU___U1338 ( .A(ALU__n1717), .Y(ALU__n1352) );
  BUFx4f_ASAP7_75t_R ALU___U1339 ( .A(ALU__N133), .Y(ALU__n1717) );
  INVx2_ASAP7_75t_R ALU___U1340 ( .A(ALU__n1723), .Y(ALU__n1331) );
  BUFx4f_ASAP7_75t_R ALU___U1341 ( .A(ALU__N127), .Y(ALU__n1723) );
  BUFx12f_ASAP7_75t_R ALU___U1342 ( .A(ALU__n715), .Y(ALU__n1449) );
  BUFx12f_ASAP7_75t_R ALU___U1343 ( .A(ALU__n860), .Y(ALU__n1642) );
  INVx3_ASAP7_75t_R ALU___U1344 ( .A(ALU__n1642), .Y(ALU__n1634) );
  CKINVDCx6p67_ASAP7_75t_R ALU___U1345 ( .A(ALU__n2), .Y(ALU__n1479) );
  INVx2_ASAP7_75t_R ALU___U1346 ( .A(ALU__n1701), .Y(ALU__n1348) );
  OR4x1_ASAP7_75t_R ALU___U1347 ( .A(EX_ALU_result[5]), .B(EX_ALU_result[4]), .C(
        EX_ALU_result[3]), .D(EX_ALU_result[31]), .Y(ALU__n124) );
  INVxp67_ASAP7_75t_R ALU___U1348 ( .A(ALU__n791), .Y(ALU__n1111) );
  BUFx2_ASAP7_75t_R ALU___U1349 ( .A(ALU__N376), .Y(ALU__n1112) );
  BUFx2_ASAP7_75t_R ALU___U1350 ( .A(ALU__n202), .Y(ALU__n1113) );
  OA221x2_ASAP7_75t_R ALU___U1351 ( .A1(ALU__n1292), .A2(ALU__n1622), .B1(ALU__n1418), .B2(ALU__n1599), 
        .C(ALU__n1234), .Y(ALU__n203) );
  INVx1_ASAP7_75t_R ALU___U1352 ( .A(ALU__n1010), .Y(ALU__n1114) );
  OA22x2_ASAP7_75t_R ALU___U1353 ( .A1(ALU__n805), .A2(ALU__n1690), .B1(n701), 
        .B2(ALU__n513), .Y(ALU__n201) );
  INVx1_ASAP7_75t_R ALU___U1354 ( .A(ALU__n1012), .Y(ALU__n1115) );
  BUFx2_ASAP7_75t_R ALU___U1355 ( .A(ALU__N369), .Y(ALU__n1116) );
  BUFx2_ASAP7_75t_R ALU___U1356 ( .A(ALU__n244), .Y(ALU__n1117) );
  OA221x2_ASAP7_75t_R ALU___U1357 ( .A1(ALU__n1378), .A2(ALU__n1620), .B1(ALU__n1014), .B2(ALU__n1601), 
        .C(ALU__n1082), .Y(ALU__n245) );
  INVx1_ASAP7_75t_R ALU___U1358 ( .A(ALU__n875), .Y(ALU__n1118) );
  OA22x2_ASAP7_75t_R ALU___U1359 ( .A1(ALU__n918), .A2(ALU__n1738), .B1(n767), 
        .B2(ALU__n580), .Y(ALU__n243) );
  INVx1_ASAP7_75t_R ALU___U1360 ( .A(ALU__n877), .Y(ALU__n1119) );
  AND4x2_ASAP7_75t_R ALU___U1361 ( .A(ALU__n1349), .B(ALU_ctl[1]), .C(ALU__n1733), .D(
        n1406), .Y(ALU__n129) );
  INVx3_ASAP7_75t_R ALU___U1362 ( .A(n794), .Y(ALU__n1697) );
  AO22x1_ASAP7_75t_R ALU___U1363 ( .A1(ALU__N166), .A2(ALU__n1562), .B1(ALU__N275), .B2(ALU__n1532), .Y(
        n228) );
  INVx2_ASAP7_75t_R ALU___U1364 ( .A(ALU__n456), .Y(ALU__n1120) );
  INVx2_ASAP7_75t_R ALU___U1365 ( .A(n892), .Y(ALU__n1700) );
  BUFx4f_ASAP7_75t_R ALU___U1366 ( .A(ALU__n1706), .Y(ALU__n1121) );
  INVx4_ASAP7_75t_R ALU___U1367 ( .A(n798), .Y(ALU__n1682) );
  BUFx12f_ASAP7_75t_R ALU___U1368 ( .A(ALU__n1464), .Y(ALU__n1122) );
  BUFx12f_ASAP7_75t_R ALU___U1369 ( .A(ALU__n1464), .Y(ALU__n1123) );
  INVx2_ASAP7_75t_R ALU___U1370 ( .A(ALU__n1708), .Y(ALU__n1351) );
  INVx2_ASAP7_75t_R ALU___U1371 ( .A(ALU__n1710), .Y(ALU__n1328) );
  INVx2_ASAP7_75t_R ALU___U1372 ( .A(ALU__n1722), .Y(ALU__n1313) );
  BUFx12f_ASAP7_75t_R ALU___U1373 ( .A(ALU__n1326), .Y(ALU__n1124) );
  BUFx6f_ASAP7_75t_R ALU___U1374 ( .A(ALU__n1326), .Y(ALU__n1125) );
  INVx5_ASAP7_75t_R ALU___U1375 ( .A(ALU__n1124), .Y(ALU__n1442) );
  INVx3_ASAP7_75t_R ALU___U1376 ( .A(ALU__n1125), .Y(ALU__n1444) );
  BUFx12f_ASAP7_75t_R ALU___U1377 ( .A(ALU__n391), .Y(ALU__n1326) );
  BUFx2_ASAP7_75t_R ALU___U1378 ( .A(ALU__n123), .Y(ALU__n1126) );
  BUFx12f_ASAP7_75t_R ALU___U1379 ( .A(n352), .Y(ALU__n1698) );
  BUFx12f_ASAP7_75t_R ALU___U1380 ( .A(ALU__n1643), .Y(ALU__n1127) );
  BUFx12f_ASAP7_75t_R ALU___U1381 ( .A(ALU__n985), .Y(ALU__n1128) );
  BUFx12f_ASAP7_75t_R ALU___U1382 ( .A(ALU__n861), .Y(ALU__n1640) );
  BUFx12f_ASAP7_75t_R ALU___U1383 ( .A(ALU__n1127), .Y(ALU__n1391) );
  BUFx12f_ASAP7_75t_R ALU___U1384 ( .A(ALU__n1644), .Y(ALU__n1643) );
  CKINVDCx8_ASAP7_75t_R ALU___U1385 ( .A(ALU__n1481), .Y(ALU__n1129) );
  BUFx12f_ASAP7_75t_R ALU___U1386 ( .A(ALU__n1497), .Y(ALU__n1130) );
  BUFx12f_ASAP7_75t_R ALU___U1387 ( .A(ALU__n47), .Y(ALU__n1497) );
  AO22x2_ASAP7_75t_R ALU___U1388 ( .A1(ALU__N164), .A2(ALU__n1561), .B1(ALU__N273), .B2(ALU__n1531), .Y(
        n240) );
  BUFx2_ASAP7_75t_R ALU___U1389 ( .A(ALU__N379), .Y(ALU__n1133) );
  BUFx2_ASAP7_75t_R ALU___U1390 ( .A(ALU__n184), .Y(ALU__n1134) );
  OA221x2_ASAP7_75t_R ALU___U1391 ( .A1(ALU__n1311), .A2(ALU__n1621), .B1(ALU__n1359), .B2(ALU__n1598), 
        .C(ALU__n605), .Y(ALU__n185) );
  INVx1_ASAP7_75t_R ALU___U1392 ( .A(ALU__n444), .Y(ALU__n1135) );
  OA22x2_ASAP7_75t_R ALU___U1393 ( .A1(ALU__n872), .A2(ALU__n1689), .B1(n1056), 
        .B2(ALU__n787), .Y(ALU__n183) );
  INVx1_ASAP7_75t_R ALU___U1394 ( .A(ALU__n446), .Y(ALU__n1136) );
  BUFx2_ASAP7_75t_R ALU___U1395 ( .A(ALU__N367), .Y(ALU__n1137) );
  BUFx2_ASAP7_75t_R ALU___U1396 ( .A(ALU__n256), .Y(ALU__n1138) );
  OA221x2_ASAP7_75t_R ALU___U1397 ( .A1(ALU__n1317), .A2(ALU__n1619), .B1(ALU__n1753), .B2(ALU__n1602), 
        .C(ALU__n958), .Y(ALU__n257) );
  INVx1_ASAP7_75t_R ALU___U1398 ( .A(ALU__n594), .Y(ALU__n1139) );
  OA22x2_ASAP7_75t_R ALU___U1399 ( .A1(ALU__n874), .A2(ALU__n1297), .B1(ALU__n80), .B2(ALU__n788), .Y(
        n255) );
  INVx1_ASAP7_75t_R ALU___U1400 ( .A(ALU__n596), .Y(ALU__n1140) );
  BUFx2_ASAP7_75t_R ALU___U1401 ( .A(ALU__N359), .Y(ALU__n1141) );
  BUFx2_ASAP7_75t_R ALU___U1402 ( .A(ALU__n304), .Y(ALU__n1142) );
  OA221x2_ASAP7_75t_R ALU___U1403 ( .A1(ALU__n1354), .A2(ALU__n1620), .B1(ALU__n1421), .B2(ALU__n1605), 
        .C(ALU__n960), .Y(ALU__n305) );
  INVx1_ASAP7_75t_R ALU___U1404 ( .A(ALU__n559), .Y(ALU__n1143) );
  OA22x2_ASAP7_75t_R ALU___U1405 ( .A1(ALU__n482), .A2(ALU__n1746), .B1(ALU__n901), .B2(ALU__n366), .Y(
        n303) );
  INVx1_ASAP7_75t_R ALU___U1406 ( .A(ALU__n561), .Y(ALU__n1144) );
  BUFx2_ASAP7_75t_R ALU___U1407 ( .A(ALU__N365), .Y(ALU__n1145) );
  BUFx2_ASAP7_75t_R ALU___U1408 ( .A(ALU__n268), .Y(ALU__n1146) );
  OA221x2_ASAP7_75t_R ALU___U1409 ( .A1(ALU__n1331), .A2(ALU__n1618), .B1(ALU__n1389), .B2(ALU__n1603), 
        .C(ALU__n1217), .Y(ALU__n269) );
  INVx1_ASAP7_75t_R ALU___U1410 ( .A(ALU__n879), .Y(ALU__n1147) );
  OA22x2_ASAP7_75t_R ALU___U1411 ( .A1(ALU__n980), .A2(ALU__n903), .B1(n1208), .B2(
        n532), .Y(ALU__n267) );
  INVx1_ASAP7_75t_R ALU___U1412 ( .A(ALU__n881), .Y(ALU__n1148) );
  AO22x2_ASAP7_75t_R ALU___U1413 ( .A1(ALU__N308), .A2(ALU__n1517), .B1(ALU__N340), .B2(ALU__n1503), .Y(
        n220) );
  BUFx2_ASAP7_75t_R ALU___U1414 ( .A(ALU__n1794), .Y(ALU__n1149) );
  BUFx2_ASAP7_75t_R ALU___U1415 ( .A(ALU__n1800), .Y(ALU__n1150) );
  BUFx2_ASAP7_75t_R ALU___U1416 ( .A(ALU__n1811), .Y(ALU__n1151) );
  AO22x2_ASAP7_75t_R ALU___U1417 ( .A1(ALU__N312), .A2(ALU__n1517), .B1(ALU__N344), .B2(ALU__n1504), .Y(
        n196) );
  BUFx12f_ASAP7_75t_R ALU___U1418 ( .A(ALU__n1154), .Y(ALU__n1152) );
  BUFx12f_ASAP7_75t_R ALU___U1419 ( .A(ALU__n1154), .Y(ALU__n1153) );
  BUFx12f_ASAP7_75t_R ALU___U1420 ( .A(ALU__n1450), .Y(ALU__n1154) );
  CKINVDCx5p33_ASAP7_75t_R ALU___U1421 ( .A(ALU__n1153), .Y(ALU__n1445) );
  CKINVDCx5p33_ASAP7_75t_R ALU___U1422 ( .A(ALU__n1152), .Y(ALU__n1434) );
  BUFx12f_ASAP7_75t_R ALU___U1423 ( .A(ALU__n1201), .Y(ALU__n1450) );
  BUFx12f_ASAP7_75t_R ALU___U1424 ( .A(ALU__n629), .Y(ALU__n1692) );
  BUFx3_ASAP7_75t_R ALU___U1425 ( .A(ALU__n1156), .Y(EX_ALU_result[10]) );
  BUFx2_ASAP7_75t_R ALU___U1426 ( .A(ALU__n1804), .Y(ALU__n1156) );
  BUFx4f_ASAP7_75t_R ALU___U1427 ( .A(ALU__n1158), .Y(EX_ALU_result[30]) );
  BUFx3_ASAP7_75t_R ALU___U1428 ( .A(ALU__n1006), .Y(ALU__n1158) );
  BUFx4f_ASAP7_75t_R ALU___U1429 ( .A(ALU__n1160), .Y(EX_ALU_result[9]) );
  BUFx3_ASAP7_75t_R ALU___U1430 ( .A(ALU__n939), .Y(ALU__n1160) );
  BUFx6f_ASAP7_75t_R ALU___U1431 ( .A(ALU__n639), .Y(ALU__n1161) );
  BUFx3_ASAP7_75t_R ALU___U1432 ( .A(ALU__n640), .Y(ALU__n1162) );
  BUFx12f_ASAP7_75t_R ALU___U1433 ( .A(ALU__n1165), .Y(ALU__n1163) );
  BUFx12f_ASAP7_75t_R ALU___U1434 ( .A(ALU__n1163), .Y(ALU__n1164) );
  BUFx12f_ASAP7_75t_R ALU___U1435 ( .A(ALU__n1468), .Y(ALU__n1165) );
  OR4x1_ASAP7_75t_R ALU___U1436 ( .A(ALU__n1406), .B(ALU__n1733), .C(ALU_ctl[1]), .D(
        ALU_ctl[0]), .Y(ALU__n139) );
  BUFx12f_ASAP7_75t_R ALU___U1437 ( .A(ALU__n1161), .Y(ALU__n1468) );
  CKINVDCx8_ASAP7_75t_R ALU___U1438 ( .A(ALU__n1536), .Y(ALU__n1167) );
  BUFx12f_ASAP7_75t_R ALU___U1439 ( .A(ALU__n1169), .Y(EX_ALU_result[27]) );
  BUFx12f_ASAP7_75t_R ALU___U1440 ( .A(ALU__n1079), .Y(ALU__n1169) );
  INVx1_ASAP7_75t_R ALU___U1441 ( .A(ALU__n474), .Y(ALU__n1170) );
  BUFx2_ASAP7_75t_R ALU___U1442 ( .A(ALU__n323), .Y(ALU__n1171) );
  BUFx2_ASAP7_75t_R ALU___U1443 ( .A(ALU__n322), .Y(ALU__n1172) );
  AO22x1_ASAP7_75t_R ALU___U1444 ( .A1(ALU__N323), .A2(ALU__n1502), .B1(ALU__N291), .B2(ALU__n1514), .Y(
        n321) );
  INVx1_ASAP7_75t_R ALU___U1445 ( .A(ALU__n476), .Y(ALU__n1173) );
  BUFx12f_ASAP7_75t_R ALU___U1446 ( .A(ALU__n63), .Y(ALU__n1174) );
  BUFx12f_ASAP7_75t_R ALU___U1447 ( .A(ALU__n64), .Y(ALU__n1175) );
  INVx6_ASAP7_75t_R ALU___U1448 ( .A(ALU__n1174), .Y(ALU__n1486) );
  BUFx3_ASAP7_75t_R ALU___U1449 ( .A(ALU__N144), .Y(ALU__n1706) );
  INVx2_ASAP7_75t_R ALU___U1450 ( .A(ALU__n1121), .Y(ALU__n1176) );
  BUFx2_ASAP7_75t_R ALU___U1451 ( .A(ALU__N380), .Y(ALU__n1177) );
  BUFx2_ASAP7_75t_R ALU___U1452 ( .A(ALU__n178), .Y(ALU__n1178) );
  OA221x2_ASAP7_75t_R ALU___U1453 ( .A1(ALU__n1351), .A2(ALU__n1621), .B1(ALU__n1392), .B2(ALU__n1598), 
        .C(ALU__n898), .Y(ALU__n179) );
  INVx1_ASAP7_75t_R ALU___U1454 ( .A(ALU__n975), .Y(ALU__n1179) );
  OA22x2_ASAP7_75t_R ALU___U1455 ( .A1(ALU__n563), .A2(ALU__n1742), .B1(n955), 
        .B2(ALU__n512), .Y(ALU__n177) );
  INVx1_ASAP7_75t_R ALU___U1456 ( .A(ALU__n977), .Y(ALU__n1180) );
  BUFx2_ASAP7_75t_R ALU___U1457 ( .A(ALU__N371), .Y(ALU__n1181) );
  BUFx2_ASAP7_75t_R ALU___U1458 ( .A(ALU__n232), .Y(ALU__n1182) );
  OA221x2_ASAP7_75t_R ALU___U1459 ( .A1(ALU__n1352), .A2(ALU__n1620), .B1(ALU__n1336), .B2(ALU__n1601), 
        .C(ALU__n1025), .Y(ALU__n233) );
  INVx1_ASAP7_75t_R ALU___U1460 ( .A(ALU__n797), .Y(ALU__n1183) );
  OA22x2_ASAP7_75t_R ALU___U1461 ( .A1(ALU__n974), .A2(ALU__n1740), .B1(n1222), 
        .B2(ALU__n818), .Y(ALU__n231) );
  INVx1_ASAP7_75t_R ALU___U1462 ( .A(ALU__n799), .Y(ALU__n1184) );
  AO22x2_ASAP7_75t_R ALU___U1463 ( .A1(ALU__N306), .A2(ALU__n1516), .B1(ALU__N338), .B2(ALU__n1504), .Y(
        n232) );
  BUFx2_ASAP7_75t_R ALU___U1464 ( .A(ALU__N363), .Y(ALU__n1185) );
  BUFx2_ASAP7_75t_R ALU___U1465 ( .A(ALU__n280), .Y(ALU__n1186) );
  OA221x2_ASAP7_75t_R ALU___U1466 ( .A1(ALU__n1315), .A2(ALU__n1618), .B1(ALU__n1275), .B2(ALU__n1603), 
        .C(ALU__n1334), .Y(ALU__n281) );
  INVx1_ASAP7_75t_R ALU___U1467 ( .A(ALU__n452), .Y(ALU__n1187) );
  OA22x2_ASAP7_75t_R ALU___U1468 ( .A1(ALU__n944), .A2(ALU__n1235), .B1(ALU__n368), .B2(ALU__n789), .Y(
        n279) );
  INVx1_ASAP7_75t_R ALU___U1469 ( .A(ALU__n454), .Y(ALU__n1188) );
  BUFx2_ASAP7_75t_R ALU___U1470 ( .A(ALU__N387), .Y(ALU__n1189) );
  BUFx2_ASAP7_75t_R ALU___U1471 ( .A(ALU__n127), .Y(ALU__n1190) );
  OA221x2_ASAP7_75t_R ALU___U1472 ( .A1(ALU__n1348), .A2(ALU__n85), .B1(ALU__n1605), .B2(ALU__n1775), 
        .C(ALU__n1038), .Y(ALU__n128) );
  INVx1_ASAP7_75t_R ALU___U1473 ( .A(ALU__n520), .Y(ALU__n1191) );
  OA22x2_ASAP7_75t_R ALU___U1474 ( .A1(ALU__n887), .A2(ALU__n1308), .B1(n888), 
        .B2(ALU__n926), .Y(ALU__n126) );
  INVx1_ASAP7_75t_R ALU___U1475 ( .A(ALU__n522), .Y(ALU__n1192) );
  INVx4_ASAP7_75t_R ALU___U1476 ( .A(n767), .Y(ALU__n1738) );
  INVx2_ASAP7_75t_R ALU___U1477 ( .A(n858), .Y(ALU__n1693) );
  CKINVDCx9p33_ASAP7_75t_R ALU___U1478 ( .A(ALU__n855), .Y(ALU__n1193) );
  BUFx12f_ASAP7_75t_R ALU___U1479 ( .A(ALU__n1193), .Y(ALU__n1586) );
  INVx4_ASAP7_75t_R ALU___U1480 ( .A(ALU__n1681), .Y(ALU__n1194) );
  BUFx2_ASAP7_75t_R ALU___U1481 ( .A(ALU__n200), .Y(ALU__n1195) );
  BUFx2_ASAP7_75t_R ALU___U1482 ( .A(ALU__n1801), .Y(ALU__n1196) );
  BUFx2_ASAP7_75t_R ALU___U1483 ( .A(ALU__n320), .Y(ALU__n1197) );
  BUFx12f_ASAP7_75t_R ALU___U1484 ( .A(ALU__n1776), .Y(ALU__n1199) );
  BUFx12f_ASAP7_75t_R ALU___U1485 ( .A(ALU__n1699), .Y(ALU__n1200) );
  BUFx12f_ASAP7_75t_R ALU___U1486 ( .A(ALU__n1203), .Y(ALU__n1201) );
  BUFx12f_ASAP7_75t_R ALU___U1487 ( .A(ALU__n1452), .Y(ALU__n1202) );
  BUFx12f_ASAP7_75t_R ALU___U1488 ( .A(ALU__n1452), .Y(ALU__n1203) );
  BUFx12f_ASAP7_75t_R ALU___U1489 ( .A(ALU__n1018), .Y(ALU__n1452) );
  BUFx3_ASAP7_75t_R ALU___U1490 ( .A(ALU__n1205), .Y(EX_ALU_result[18]) );
  BUFx2_ASAP7_75t_R ALU___U1491 ( .A(ALU__n1796), .Y(ALU__n1205) );
  BUFx4f_ASAP7_75t_R ALU___U1492 ( .A(ALU__n1209), .Y(EX_ALU_result[29]) );
  BUFx3_ASAP7_75t_R ALU___U1493 ( .A(ALU__n1068), .Y(ALU__n1209) );
  BUFx4f_ASAP7_75t_R ALU___U1494 ( .A(ALU__n1211), .Y(EX_ALU_result[22]) );
  BUFx3_ASAP7_75t_R ALU___U1495 ( .A(ALU__n841), .Y(ALU__n1211) );
  BUFx4f_ASAP7_75t_R ALU___U1496 ( .A(ALU__n1213), .Y(EX_ALU_result[6]) );
  BUFx3_ASAP7_75t_R ALU___U1497 ( .A(ALU__n1045), .Y(ALU__n1213) );
  BUFx12f_ASAP7_75t_R ALU___U1498 ( .A(ALU__n1215), .Y(EX_ALU_result[25]) );
  BUFx12f_ASAP7_75t_R ALU___U1499 ( .A(ALU__n1058), .Y(ALU__n1215) );
  INVx3_ASAP7_75t_R ALU___U1500 ( .A(ALU__n1696), .Y(ALU__n1216) );
  AO22x1_ASAP7_75t_R ALU___U1501 ( .A1(ALU__N159), .A2(ALU__n1559), .B1(ALU__N268), .B2(ALU__n1529), .Y(
        n270) );
  BUFx2_ASAP7_75t_R ALU___U1502 ( .A(ALU__N366), .Y(ALU__n1218) );
  BUFx2_ASAP7_75t_R ALU___U1503 ( .A(ALU__n262), .Y(ALU__n1219) );
  OA221x2_ASAP7_75t_R ALU___U1504 ( .A1(ALU__n1313), .A2(ALU__n1619), .B1(ALU__n1386), .B2(ALU__n1601), 
        .C(ALU__n989), .Y(ALU__n263) );
  INVx1_ASAP7_75t_R ALU___U1505 ( .A(ALU__n949), .Y(ALU__n1220) );
  OA22x2_ASAP7_75t_R ALU___U1506 ( .A1(ALU__n919), .A2(ALU__n1005), .B1(n1164), 
        .B2(ALU__n433), .Y(ALU__n261) );
  INVx1_ASAP7_75t_R ALU___U1507 ( .A(ALU__n951), .Y(ALU__n1221) );
  BUFx2_ASAP7_75t_R ALU___U1508 ( .A(ALU__N360), .Y(ALU__n1222) );
  BUFx2_ASAP7_75t_R ALU___U1509 ( .A(ALU__n298), .Y(ALU__n1223) );
  OA221x2_ASAP7_75t_R ALU___U1510 ( .A1(ALU__n1332), .A2(ALU__n1618), .B1(ALU__n1360), .B2(ALU__n1604), 
        .C(ALU__n706), .Y(ALU__n299) );
  INVx1_ASAP7_75t_R ALU___U1511 ( .A(ALU__n478), .Y(ALU__n1224) );
  OA22x2_ASAP7_75t_R ALU___U1512 ( .A1(ALU__n1307), .A2(ALU__n1747), .B1(ALU__n783), .B2(ALU__n790), .Y(
        n297) );
  INVx1_ASAP7_75t_R ALU___U1513 ( .A(ALU__n480), .Y(ALU__n1225) );
  BUFx2_ASAP7_75t_R ALU___U1514 ( .A(ALU__N384), .Y(ALU__n1226) );
  OA221x2_ASAP7_75t_R ALU___U1515 ( .A1(ALU__n1704), .A2(ALU__n1623), .B1(ALU__n1420), .B2(ALU__n1597), 
        .C(ALU__n990), .Y(ALU__n155) );
  INVx1_ASAP7_75t_R ALU___U1516 ( .A(ALU__n551), .Y(ALU__n1227) );
  BUFx2_ASAP7_75t_R ALU___U1517 ( .A(ALU__n154), .Y(ALU__n1228) );
  OA22x2_ASAP7_75t_R ALU___U1518 ( .A1(ALU__n1306), .A2(ALU__n1105), .B1(n1033), 
        .B2(ALU__n1008), .Y(ALU__n153) );
  INVx1_ASAP7_75t_R ALU___U1519 ( .A(ALU__n553), .Y(ALU__n1229) );
  INVx2_ASAP7_75t_R ALU___U1520 ( .A(ALU__N146), .Y(ALU__n1704) );
  BUFx2_ASAP7_75t_R ALU___U1521 ( .A(ALU__N382), .Y(ALU__n1230) );
  BUFx2_ASAP7_75t_R ALU___U1522 ( .A(ALU__n166), .Y(ALU__n1231) );
  OA221x2_ASAP7_75t_R ALU___U1523 ( .A1(ALU__n1176), .A2(ALU__n1622), .B1(ALU__n1419), .B2(ALU__n1598), 
        .C(ALU__n681), .Y(ALU__n167) );
  INVx1_ASAP7_75t_R ALU___U1524 ( .A(ALU__n421), .Y(ALU__n1232) );
  OA22x2_ASAP7_75t_R ALU___U1525 ( .A1(ALU__n925), .A2(ALU__n1066), .B1(n978), 
        .B2(ALU__n814), .Y(ALU__n165) );
  INVx1_ASAP7_75t_R ALU___U1526 ( .A(ALU__n423), .Y(ALU__n1233) );
  AO22x1_ASAP7_75t_R ALU___U1527 ( .A1(ALU__N170), .A2(ALU__n1563), .B1(ALU__N279), .B2(ALU__n1528), .Y(
        n204) );
  INVx4_ASAP7_75t_R ALU___U1528 ( .A(ALU__n1748), .Y(ALU__n1235) );
  AO22x2_ASAP7_75t_R ALU___U1529 ( .A1(ALU__N309), .A2(ALU__n1517), .B1(ALU__N341), .B2(ALU__n1504), .Y(
        n214) );
  BUFx6f_ASAP7_75t_R ALU___U1530 ( .A(ALU__n1466), .Y(ALU__n1455) );
  BUFx4f_ASAP7_75t_R ALU___U1531 ( .A(ALU__n1030), .Y(ALU__n1773) );
  BUFx12f_ASAP7_75t_R ALU___U1532 ( .A(ALU__n1769), .Y(ALU__n1236) );
  BUFx12f_ASAP7_75t_R ALU___U1533 ( .A(ALU__n1756), .Y(ALU__n1237) );
  BUFx12f_ASAP7_75t_R ALU___U1534 ( .A(ALU__n1782), .Y(ALU__n1238) );
  BUFx3_ASAP7_75t_R ALU___U1535 ( .A(ALU__n1242), .Y(EX_ALU_result[0]) );
  BUFx2_ASAP7_75t_R ALU___U1536 ( .A(ALU__n1814), .Y(ALU__n1242) );
  BUFx4f_ASAP7_75t_R ALU___U1537 ( .A(ALU__n1244), .Y(EX_ALU_result[28]) );
  BUFx3_ASAP7_75t_R ALU___U1538 ( .A(ALU__n840), .Y(ALU__n1244) );
  BUFx4f_ASAP7_75t_R ALU___U1539 ( .A(ALU__n1246), .Y(EX_ALU_result[23]) );
  BUFx3_ASAP7_75t_R ALU___U1540 ( .A(ALU__n1044), .Y(ALU__n1246) );
  BUFx4f_ASAP7_75t_R ALU___U1541 ( .A(ALU__n1248), .Y(EX_ALU_result[15]) );
  BUFx3_ASAP7_75t_R ALU___U1542 ( .A(ALU__n1070), .Y(ALU__n1248) );
  BUFx4f_ASAP7_75t_R ALU___U1543 ( .A(ALU__n1250), .Y(EX_ALU_result[8]) );
  BUFx3_ASAP7_75t_R ALU___U1544 ( .A(ALU__n1007), .Y(ALU__n1250) );
  BUFx12f_ASAP7_75t_R ALU___U1545 ( .A(ALU__n1790), .Y(EX_ALU_result[24]) );
  INVx4_ASAP7_75t_R ALU___U1546 ( .A(n1075), .Y(ALU__n1741) );
  INVx4_ASAP7_75t_R ALU___U1547 ( .A(ALU__n899), .Y(ALU__n1746) );
  BUFx2_ASAP7_75t_R ALU___U1548 ( .A(ALU__N119), .Y(ALU__n1731) );
  INVx1_ASAP7_75t_R ALU___U1549 ( .A(ALU__n1731), .Y(ALU__n1253) );
  BUFx12f_ASAP7_75t_R ALU___U1550 ( .A(ALU__n1257), .Y(ALU__n1255) );
  BUFx12f_ASAP7_75t_R ALU___U1551 ( .A(ALU__n1498), .Y(ALU__n1257) );
  BUFx12f_ASAP7_75t_R ALU___U1552 ( .A(ALU__n1498), .Y(ALU__n1258) );
  BUFx12f_ASAP7_75t_R ALU___U1553 ( .A(ALU__n1395), .Y(ALU__n1498) );
  BUFx2_ASAP7_75t_R ALU___U1554 ( .A(ALU__N378), .Y(ALU__n1259) );
  BUFx2_ASAP7_75t_R ALU___U1555 ( .A(ALU__n190), .Y(ALU__n1260) );
  OA221x2_ASAP7_75t_R ALU___U1556 ( .A1(ALU__n1328), .A2(ALU__n1621), .B1(ALU__n1393), .B2(ALU__n1597), 
        .C(ALU__n707), .Y(ALU__n191) );
  INVx1_ASAP7_75t_R ALU___U1557 ( .A(ALU__n434), .Y(ALU__n1261) );
  OA22x2_ASAP7_75t_R ALU___U1558 ( .A1(ALU__n953), .A2(ALU__n1106), .B1(n1162), 
        .B2(ALU__n473), .Y(ALU__n189) );
  INVx1_ASAP7_75t_R ALU___U1559 ( .A(ALU__n436), .Y(ALU__n1262) );
  BUFx2_ASAP7_75t_R ALU___U1560 ( .A(ALU__N372), .Y(ALU__n1263) );
  OA221x2_ASAP7_75t_R ALU___U1561 ( .A1(ALU__n1716), .A2(ALU__n1622), .B1(ALU__n981), .B2(ALU__n1600), 
        .C(ALU__n1120), .Y(ALU__n227) );
  INVx1_ASAP7_75t_R ALU___U1562 ( .A(ALU__n535), .Y(ALU__n1264) );
  BUFx2_ASAP7_75t_R ALU___U1563 ( .A(ALU__n226), .Y(ALU__n1265) );
  OA22x2_ASAP7_75t_R ALU___U1564 ( .A1(ALU__n943), .A2(ALU__n1695), .B1(n547), 
        .B2(ALU__n866), .Y(ALU__n225) );
  INVx1_ASAP7_75t_R ALU___U1565 ( .A(ALU__n537), .Y(ALU__n1266) );
  INVx2_ASAP7_75t_R ALU___U1566 ( .A(ALU__N134), .Y(ALU__n1716) );
  INVx4_ASAP7_75t_R ALU___U1567 ( .A(n547), .Y(ALU__n1695) );
  BUFx2_ASAP7_75t_R ALU___U1568 ( .A(ALU__N361), .Y(ALU__n1267) );
  BUFx2_ASAP7_75t_R ALU___U1569 ( .A(ALU__n292), .Y(ALU__n1268) );
  OA221x2_ASAP7_75t_R ALU___U1570 ( .A1(ALU__n1727), .A2(ALU__n1621), .B1(ALU__n1387), .B2(ALU__n1604), 
        .C(ALU__n1293), .Y(ALU__n293) );
  INVx1_ASAP7_75t_R ALU___U1571 ( .A(ALU__n827), .Y(ALU__n1269) );
  OA22x2_ASAP7_75t_R ALU___U1572 ( .A1(ALU__n920), .A2(ALU__n1682), .B1(n798), .B2(
        n864), .Y(ALU__n291) );
  INVx1_ASAP7_75t_R ALU___U1573 ( .A(ALU__n829), .Y(ALU__n1270) );
  INVx2_ASAP7_75t_R ALU___U1574 ( .A(ALU__N123), .Y(ALU__n1727) );
  CKINVDCx9p33_ASAP7_75t_R ALU___U1575 ( .A(ALU__n809), .Y(ALU__n1271) );
  BUFx12f_ASAP7_75t_R ALU___U1576 ( .A(ALU__n1274), .Y(ALU__n1272) );
  BUFx12f_ASAP7_75t_R ALU___U1577 ( .A(ALU__n839), .Y(ALU__n1273) );
  BUFx12f_ASAP7_75t_R ALU___U1578 ( .A(ALU__n1506), .Y(ALU__n1274) );
  BUFx12f_ASAP7_75t_R ALU___U1579 ( .A(ALU__n632), .Y(ALU__n1511) );
  BUFx12f_ASAP7_75t_R ALU___U1580 ( .A(ALU__n631), .Y(ALU__n1510) );
  BUFx12f_ASAP7_75t_R ALU___U1581 ( .A(ALU__n711), .Y(ALU__n1509) );
  BUFx6f_ASAP7_75t_R ALU___U1582 ( .A(n1114), .Y(ALU__n1780) );
  INVx4_ASAP7_75t_R ALU___U1583 ( .A(ALU__n749), .Y(ALU__n1275) );
  BUFx4f_ASAP7_75t_R ALU___U1584 ( .A(ALU__n1277), .Y(ALU__n1276) );
  BUFx3_ASAP7_75t_R ALU___U1585 ( .A(ALU__n606), .Y(ALU__n1277) );
  AO22x2_ASAP7_75t_R ALU___U1586 ( .A1(ALU__N310), .A2(ALU__n1517), .B1(ALU__N342), .B2(ALU__n1505), .Y(
        n208) );
  BUFx4f_ASAP7_75t_R ALU___U1587 ( .A(ALU__n1281), .Y(EX_ALU_result[21]) );
  BUFx3_ASAP7_75t_R ALU___U1588 ( .A(ALU__n1069), .Y(ALU__n1281) );
  BUFx4f_ASAP7_75t_R ALU___U1589 ( .A(ALU__n1283), .Y(EX_ALU_result[16]) );
  BUFx3_ASAP7_75t_R ALU___U1590 ( .A(ALU__n842), .Y(ALU__n1283) );
  BUFx4f_ASAP7_75t_R ALU___U1591 ( .A(ALU__n1285), .Y(EX_ALU_result[2]) );
  BUFx3_ASAP7_75t_R ALU___U1592 ( .A(ALU__n1046), .Y(ALU__n1285) );
  BUFx12f_ASAP7_75t_R ALU___U1593 ( .A(ALU__n1451), .Y(ALU__n1286) );
  BUFx12f_ASAP7_75t_R ALU___U1594 ( .A(ALU__n376), .Y(ALU__n1287) );
  CKINVDCx5p33_ASAP7_75t_R ALU___U1595 ( .A(ALU__n1286), .Y(ALU__n1433) );
  BUFx12f_ASAP7_75t_R ALU___U1596 ( .A(ALU__n760), .Y(ALU__n1451) );
  BUFx3_ASAP7_75t_R ALU___U1597 ( .A(ALU__n1691), .Y(ALU__n1288) );
  BUFx2_ASAP7_75t_R ALU___U1598 ( .A(ALU__n1691), .Y(ALU__n1289) );
  INVx2_ASAP7_75t_R ALU___U1599 ( .A(n749), .Y(ALU__n1691) );
  BUFx12f_ASAP7_75t_R ALU___U1600 ( .A(ALU__n1788), .Y(EX_ALU_result[26]) );
  OR4x1_ASAP7_75t_R ALU___U1601 ( .A(EX_ALU_result[9]), .B(EX_ALU_result[8]), .C(
        EX_ALU_result[7]), .D(EX_ALU_result[6]), .Y(ALU__n125) );
  INVxp67_ASAP7_75t_R ALU___U1602 ( .A(ALU__n819), .Y(ALU__n1291) );
  BUFx2_ASAP7_75t_R ALU___U1603 ( .A(ALU__N138), .Y(ALU__n1712) );
  CKINVDCx12_ASAP7_75t_R ALU___U1604 ( .A(ALU__n1624), .Y(ALU__n1294) );
  CKINVDCx8_ASAP7_75t_R ALU___U1605 ( .A(ALU__n1619), .Y(ALU__n1295) );
  BUFx12f_ASAP7_75t_R ALU___U1606 ( .A(ALU__n500), .Y(ALU__n1611) );
  INVx6_ASAP7_75t_R ALU___U1607 ( .A(ALU__n858), .Y(ALU__n1594) );
  INVx6_ASAP7_75t_R ALU___U1608 ( .A(ALU__n705), .Y(ALU__n1587) );
  INVx4_ASAP7_75t_R ALU___U1609 ( .A(ALU__n1200), .Y(ALU__n1297) );
  INVx4_ASAP7_75t_R ALU___U1610 ( .A(ALU__n1692), .Y(ALU__n1298) );
  OR4x2_ASAP7_75t_R ALU___U1611 ( .A(ALU__n988), .B(ALU__n1406), .C(ALU_ctl[3]), .D(
        ALU_ctl[0]), .Y(ALU__n1299) );
  BUFx12f_ASAP7_75t_R ALU___U1612 ( .A(ALU__n1761), .Y(ALU__n1300) );
  BUFx6f_ASAP7_75t_R ALU___U1613 ( .A(ALU__n1773), .Y(ALU__n1416) );
  BUFx16f_ASAP7_75t_R ALU___U1614 ( .A(ALU__n1508), .Y(ALU__n1507) );
  BUFx12f_ASAP7_75t_R ALU___U1615 ( .A(ALU__n710), .Y(ALU__n1508) );
  CKINVDCx8_ASAP7_75t_R ALU___U1616 ( .A(ALU__n1509), .Y(ALU__n1504) );
  CKINVDCx8_ASAP7_75t_R ALU___U1617 ( .A(ALU__n1510), .Y(ALU__n1503) );
  BUFx4f_ASAP7_75t_R ALU___U1618 ( .A(ALU__n1303), .Y(EX_ALU_result[20]) );
  BUFx3_ASAP7_75t_R ALU___U1619 ( .A(ALU__n1149), .Y(ALU__n1303) );
  BUFx4f_ASAP7_75t_R ALU___U1620 ( .A(ALU__n1305), .Y(EX_ALU_result[14]) );
  BUFx3_ASAP7_75t_R ALU___U1621 ( .A(ALU__n1150), .Y(ALU__n1305) );
  BUFx2_ASAP7_75t_R ALU___U1622 ( .A(ALU__n157), .Y(ALU__n1306) );
  BUFx2_ASAP7_75t_R ALU___U1623 ( .A(ALU__n301), .Y(ALU__n1307) );
  BUFx6f_ASAP7_75t_R ALU___U1624 ( .A(n888), .Y(ALU__n1745) );
  INVx3_ASAP7_75t_R ALU___U1625 ( .A(ALU__n1745), .Y(ALU__n1308) );
  AND2x2_ASAP7_75t_R ALU___U1626 ( .A(ALU__n1733), .B(ALU__n668), .Y(ALU__n327) );
  INVx2_ASAP7_75t_R ALU___U1627 ( .A(ALU__n1276), .Y(ALU__n1309) );
  BUFx2_ASAP7_75t_R ALU___U1628 ( .A(ALU__N147), .Y(ALU__n1703) );
  INVx1_ASAP7_75t_R ALU___U1629 ( .A(ALU__n1703), .Y(ALU__n1310) );
  BUFx2_ASAP7_75t_R ALU___U1630 ( .A(ALU__N141), .Y(ALU__n1709) );
  BUFx2_ASAP7_75t_R ALU___U1631 ( .A(ALU__N139), .Y(ALU__n1711) );
  INVx1_ASAP7_75t_R ALU___U1632 ( .A(ALU__n1711), .Y(ALU__n1312) );
  BUFx2_ASAP7_75t_R ALU___U1633 ( .A(ALU__N128), .Y(ALU__n1722) );
  BUFx2_ASAP7_75t_R ALU___U1634 ( .A(ALU__N130), .Y(ALU__n1720) );
  INVx1_ASAP7_75t_R ALU___U1635 ( .A(ALU__n1720), .Y(ALU__n1314) );
  BUFx2_ASAP7_75t_R ALU___U1636 ( .A(ALU__N125), .Y(ALU__n1725) );
  BUFx2_ASAP7_75t_R ALU___U1637 ( .A(ALU__N129), .Y(ALU__n1721) );
  INVx4_ASAP7_75t_R ALU___U1638 ( .A(n851), .Y(ALU__n1687) );
  BUFx2_ASAP7_75t_R ALU___U1639 ( .A(ALU__n1346), .Y(ALU__n1319) );
  AO22x2_ASAP7_75t_R ALU___U1640 ( .A1(ALU__N307), .A2(ALU__n1517), .B1(ALU__N339), .B2(ALU__n1502), .Y(
        n226) );
  BUFx12f_ASAP7_75t_R ALU___U1641 ( .A(ALU__n1781), .Y(ALU__n1320) );
  BUFx12f_ASAP7_75t_R ALU___U1642 ( .A(ALU__n1123), .Y(ALU__n1321) );
  BUFx12f_ASAP7_75t_R ALU___U1643 ( .A(ALU__n1122), .Y(ALU__n1322) );
  BUFx12f_ASAP7_75t_R ALU___U1644 ( .A(ALU__n1467), .Y(ALU__n1464) );
  BUFx4f_ASAP7_75t_R ALU___U1645 ( .A(ALU__n1324), .Y(EX_ALU_result[13]) );
  BUFx3_ASAP7_75t_R ALU___U1646 ( .A(ALU__n1196), .Y(ALU__n1324) );
  AO22x2_ASAP7_75t_R ALU___U1647 ( .A1(ALU__N321), .A2(ALU__n1519), .B1(ALU__N353), .B2(ALU__n1502), .Y(
        n142) );
  AO22x2_ASAP7_75t_R ALU___U1648 ( .A1(ALU__N318), .A2(ALU__n1518), .B1(ALU__N350), .B2(ALU__n1505), .Y(
        n160) );
  INVx4_ASAP7_75t_R ALU___U1649 ( .A(ALU__n1520), .Y(ALU__n1519) );
  BUFx12f_ASAP7_75t_R ALU___U1650 ( .A(ALU__n700), .Y(ALU__n1520) );
  BUFx12f_ASAP7_75t_R ALU___U1651 ( .A(ALU__n391), .Y(ALU__n1325) );
  BUFx12f_ASAP7_75t_R ALU___U1652 ( .A(ALU__n761), .Y(ALU__n1327) );
  BUFx2_ASAP7_75t_R ALU___U1653 ( .A(ALU__N140), .Y(ALU__n1710) );
  BUFx2_ASAP7_75t_R ALU___U1654 ( .A(ALU__N136), .Y(ALU__n1714) );
  INVx1_ASAP7_75t_R ALU___U1655 ( .A(ALU__n1714), .Y(ALU__n1329) );
  BUFx2_ASAP7_75t_R ALU___U1656 ( .A(ALU__N135), .Y(ALU__n1715) );
  INVx1_ASAP7_75t_R ALU___U1657 ( .A(ALU__n1715), .Y(ALU__n1330) );
  BUFx2_ASAP7_75t_R ALU___U1658 ( .A(ALU__N122), .Y(ALU__n1728) );
  INVx1_ASAP7_75t_R ALU___U1659 ( .A(ALU__n1728), .Y(ALU__n1332) );
  BUFx2_ASAP7_75t_R ALU___U1660 ( .A(ALU__N137), .Y(ALU__n1713) );
  INVx1_ASAP7_75t_R ALU___U1661 ( .A(ALU__n1713), .Y(ALU__n1333) );
  BUFx6f_ASAP7_75t_R ALU___U1662 ( .A(n1225), .Y(ALU__n1764) );
  BUFx5_ASAP7_75t_R ALU___U1663 ( .A(n925), .Y(ALU__n1757) );
  BUFx5_ASAP7_75t_R ALU___U1664 ( .A(n969), .Y(ALU__n1756) );
  INVx4_ASAP7_75t_R ALU___U1665 ( .A(ALU__n1500), .Y(ALU__n1478) );
  BUFx12f_ASAP7_75t_R ALU___U1666 ( .A(ALU__n1256), .Y(ALU__n1493) );
  BUFx6f_ASAP7_75t_R ALU___U1667 ( .A(ALU__n1343), .Y(ALU__n1513) );
  BUFx4f_ASAP7_75t_R ALU___U1668 ( .A(ALU__n1344), .Y(ALU__n1343) );
  BUFx3_ASAP7_75t_R ALU___U1669 ( .A(ALU__n458), .Y(ALU__n1344) );
  BUFx12f_ASAP7_75t_R ALU___U1670 ( .A(ALU__n1342), .Y(ALU__n1512) );
  INVx4_ASAP7_75t_R ALU___U1671 ( .A(ALU__n1698), .Y(ALU__n1345) );
  BUFx2_ASAP7_75t_R ALU___U1672 ( .A(ALU__n1404), .Y(ALU__n1374) );
  INVx1_ASAP7_75t_R ALU___U1673 ( .A(ALU__n1374), .Y(ALU__n1346) );
  BUFx2_ASAP7_75t_R ALU___U1674 ( .A(ALU__n117), .Y(ALU__n1347) );
  BUFx6f_ASAP7_75t_R ALU___U1675 ( .A(ALU__n1465), .Y(ALU__n1458) );
  BUFx6f_ASAP7_75t_R ALU___U1676 ( .A(ALU__n1465), .Y(ALU__n1457) );
  BUFx6f_ASAP7_75t_R ALU___U1677 ( .A(ALU__n1465), .Y(ALU__n1456) );
  BUFx12f_ASAP7_75t_R ALU___U1678 ( .A(ALU__n1040), .Y(ALU__n1465) );
  BUFx2_ASAP7_75t_R ALU___U1679 ( .A(ALU__N143), .Y(ALU__n1707) );
  INVx1_ASAP7_75t_R ALU___U1680 ( .A(ALU__n1707), .Y(ALU__n1350) );
  BUFx2_ASAP7_75t_R ALU___U1681 ( .A(ALU__N142), .Y(ALU__n1708) );
  BUFx2_ASAP7_75t_R ALU___U1682 ( .A(ALU__N132), .Y(ALU__n1718) );
  BUFx2_ASAP7_75t_R ALU___U1683 ( .A(ALU__N121), .Y(ALU__n1729) );
  BUFx2_ASAP7_75t_R ALU___U1684 ( .A(ALU__N126), .Y(ALU__n1724) );
  INVx1_ASAP7_75t_R ALU___U1685 ( .A(ALU__n1724), .Y(ALU__n1355) );
  BUFx16f_ASAP7_75t_R ALU___U1686 ( .A(ALU__n1553), .Y(ALU__n1544) );
  BUFx16f_ASAP7_75t_R ALU___U1687 ( .A(ALU__n853), .Y(ALU__n1543) );
  BUFx16f_ASAP7_75t_R ALU___U1688 ( .A(ALU__n774), .Y(ALU__n1541) );
  BUFx16f_ASAP7_75t_R ALU___U1689 ( .A(ALU__n1554), .Y(ALU__n1540) );
  BUFx12f_ASAP7_75t_R ALU___U1690 ( .A(ALU__n1167), .Y(ALU__n1554) );
  CKINVDCx8_ASAP7_75t_R ALU___U1691 ( .A(ALU__n1432), .Y(ALU__n1357) );
  INVx4_ASAP7_75t_R ALU___U1692 ( .A(ALU__n1357), .Y(ALU__n1436) );
  INVx4_ASAP7_75t_R ALU___U1693 ( .A(ALU__n1357), .Y(ALU__n1435) );
  BUFx6f_ASAP7_75t_R ALU___U1694 ( .A(n1215), .Y(ALU__n1772) );
  BUFx6f_ASAP7_75t_R ALU___U1695 ( .A(n1178), .Y(ALU__n1766) );
  BUFx6f_ASAP7_75t_R ALU___U1696 ( .A(n1174), .Y(ALU__n1777) );
  BUFx6f_ASAP7_75t_R ALU___U1697 ( .A(n1182), .Y(ALU__n1760) );
  BUFx4f_ASAP7_75t_R ALU___U1698 ( .A(n1160), .Y(ALU__n1770) );
  BUFx5_ASAP7_75t_R ALU___U1699 ( .A(n973), .Y(ALU__n1779) );
  INVx2_ASAP7_75t_R ALU___U1700 ( .A(ALU__n906), .Y(ALU__n1639) );
  INVx2_ASAP7_75t_R ALU___U1701 ( .A(ALU__n1643), .Y(ALU__n1638) );
  INVx2_ASAP7_75t_R ALU___U1702 ( .A(ALU__n1644), .Y(ALU__n1637) );
  INVx3_ASAP7_75t_R ALU___U1703 ( .A(ALU__n1391), .Y(ALU__n1635) );
  INVx3_ASAP7_75t_R ALU___U1704 ( .A(ALU__n1640), .Y(ALU__n1636) );
  BUFx12f_ASAP7_75t_R ALU___U1705 ( .A(ALU__n29), .Y(ALU__n1609) );
  BUFx12f_ASAP7_75t_R ALU___U1706 ( .A(ALU__n53), .Y(ALU__n1366) );
  BUFx12f_ASAP7_75t_R ALU___U1707 ( .A(ALU__n52), .Y(ALU__n1367) );
  BUFx12f_ASAP7_75t_R ALU___U1708 ( .A(ALU__n58), .Y(ALU__n1368) );
  BUFx12f_ASAP7_75t_R ALU___U1709 ( .A(ALU__n57), .Y(ALU__n1369) );
  BUFx12f_ASAP7_75t_R ALU___U1710 ( .A(ALU__n114), .Y(ALU__n1370) );
  BUFx12f_ASAP7_75t_R ALU___U1711 ( .A(ALU__n113), .Y(ALU__n1371) );
  INVx6_ASAP7_75t_R ALU___U1712 ( .A(ALU__n1369), .Y(ALU__n1490) );
  INVx6_ASAP7_75t_R ALU___U1713 ( .A(ALU__n1368), .Y(ALU__n1489) );
  INVx6_ASAP7_75t_R ALU___U1714 ( .A(ALU__n1367), .Y(ALU__n1488) );
  INVx6_ASAP7_75t_R ALU___U1715 ( .A(ALU__n1366), .Y(ALU__n1487) );
  BUFx12f_ASAP7_75t_R ALU___U1716 ( .A(ALU__n48), .Y(ALU__n1491) );
  INVx5_ASAP7_75t_R ALU___U1717 ( .A(ALU__n1751), .Y(ALU__n1372) );
  AND2x2_ASAP7_75t_R ALU___U1718 ( .A(ALU__n1402), .B(ALU__n1403), .Y(ALU__n117) );
  INVx1_ASAP7_75t_R ALU___U1719 ( .A(ALU__n1347), .Y(ALU__n1373) );
  AND2x2_ASAP7_75t_R ALU___U1720 ( .A(ALU__n867), .B(ALU__n1410), .Y(ALU__n1404) );
  BUFx2_ASAP7_75t_R ALU___U1721 ( .A(ALU__n1405), .Y(ALU__n1375) );
  INVx1_ASAP7_75t_R ALU___U1722 ( .A(ALU__n1319), .Y(ALU__n1402) );
  INVx1_ASAP7_75t_R ALU___U1723 ( .A(ALU__n1375), .Y(ALU__n1403) );
  NAND2xp33_ASAP7_75t_R ALU___U1724 ( .A(ALU__n1111), .B(ALU__n1291), .Y(ALU__n1405) );
  BUFx12f_ASAP7_75t_R ALU___U1725 ( .A(ALU__n1762), .Y(ALU__n1376) );
  BUFx12f_ASAP7_75t_R ALU___U1726 ( .A(ALU__n1101), .Y(ALU__n1466) );
  BUFx12f_ASAP7_75t_R ALU___U1727 ( .A(ALU__n1164), .Y(ALU__n1467) );
  AO22x2_ASAP7_75t_R ALU___U1728 ( .A1(ALU__N319), .A2(ALU__n1519), .B1(ALU__N351), .B2(ALU__n1503), .Y(
        n154) );
  BUFx2_ASAP7_75t_R ALU___U1729 ( .A(ALU__N120), .Y(ALU__n1730) );
  INVx1_ASAP7_75t_R ALU___U1730 ( .A(ALU__n1730), .Y(ALU__n1377) );
  BUFx2_ASAP7_75t_R ALU___U1731 ( .A(ALU__N131), .Y(ALU__n1719) );
  INVx1_ASAP7_75t_R ALU___U1732 ( .A(ALU__n1719), .Y(ALU__n1378) );
  BUFx16f_ASAP7_75t_R ALU___U1733 ( .A(ALU__n1380), .Y(ALU__n1574) );
  BUFx16f_ASAP7_75t_R ALU___U1734 ( .A(ALU__n775), .Y(ALU__n1572) );
  BUFx12f_ASAP7_75t_R ALU___U1735 ( .A(ALU__n1581), .Y(ALU__n1585) );
  BUFx4f_ASAP7_75t_R ALU___U1736 ( .A(ALU__n1382), .Y(EX_ALU_result[7]) );
  BUFx3_ASAP7_75t_R ALU___U1737 ( .A(ALU__n1071), .Y(ALU__n1382) );
  BUFx4f_ASAP7_75t_R ALU___U1738 ( .A(ALU__n1384), .Y(EX_ALU_result[3]) );
  BUFx3_ASAP7_75t_R ALU___U1739 ( .A(ALU__n1151), .Y(ALU__n1384) );
  BUFx6f_ASAP7_75t_R ALU___U1740 ( .A(n1229), .Y(ALU__n1752) );
  BUFx6f_ASAP7_75t_R ALU___U1741 ( .A(n1233), .Y(ALU__n1778) );
  BUFx6f_ASAP7_75t_R ALU___U1742 ( .A(ALU__n965), .Y(ALU__n1759) );
  INVx4_ASAP7_75t_R ALU___U1743 ( .A(ALU__n1759), .Y(ALU__n1388) );
  BUFx5_ASAP7_75t_R ALU___U1744 ( .A(n1029), .Y(ALU__n1782) );
  BUFx5_ASAP7_75t_R ALU___U1745 ( .A(n929), .Y(ALU__n1781) );
  INVx3_ASAP7_75t_R ALU___U1746 ( .A(ALU__n779), .Y(ALU__n1596) );
  BUFx12f_ASAP7_75t_R ALU___U1747 ( .A(ALU__n28), .Y(ALU__n1608) );
  INVx4_ASAP7_75t_R ALU___U1748 ( .A(ALU__n333), .Y(ALU__n1438) );
  INVx4_ASAP7_75t_R ALU___U1749 ( .A(ALU__n332), .Y(ALU__n1437) );
  BUFx12f_ASAP7_75t_R ALU___U1750 ( .A(ALU__n1449), .Y(ALU__n1448) );
  INVx6_ASAP7_75t_R ALU___U1751 ( .A(ALU__n1325), .Y(ALU__n1443) );
  INVx2_ASAP7_75t_R ALU___U1752 ( .A(ALU__n1127), .Y(ALU__n1632) );
  INVx2_ASAP7_75t_R ALU___U1753 ( .A(ALU__n1391), .Y(ALU__n1631) );
  INVx2_ASAP7_75t_R ALU___U1754 ( .A(ALU__n861), .Y(ALU__n1630) );
  INVx2_ASAP7_75t_R ALU___U1755 ( .A(ALU__n1642), .Y(ALU__n1629) );
  INVx2_ASAP7_75t_R ALU___U1756 ( .A(ALU__n1640), .Y(ALU__n1628) );
  BUFx5_ASAP7_75t_R ALU___U1757 ( .A(n1064), .Y(ALU__n1767) );
  BUFx5_ASAP7_75t_R ALU___U1758 ( .A(n1024), .Y(ALU__n1765) );
  INVx5_ASAP7_75t_R ALU___U1759 ( .A(ALU__n1470), .Y(ALU__n1395) );
  BUFx6f_ASAP7_75t_R ALU___U1760 ( .A(ALU__n338), .Y(ALU__n1501) );
  INVx2_ASAP7_75t_R ALU___U1761 ( .A(ALU__n698), .Y(ALU__n1397) );
  BUFx12f_ASAP7_75t_R ALU___U1762 ( .A(ALU__n1396), .Y(ALU__n1500) );
  BUFx12f_ASAP7_75t_R ALU___U1763 ( .A(ALU__n1500), .Y(ALU__n1499) );
  BUFx2_ASAP7_75t_R ALU___U1764 ( .A(ALU__n118), .Y(ALU__n1400) );
  BUFx2_ASAP7_75t_R ALU___U1765 ( .A(ALU__n119), .Y(ALU__n1401) );
  OR4x1_ASAP7_75t_R ALU___U1766 ( .A(EX_ALU_result[30]), .B(EX_ALU_result[2]), .C(
        EX_ALU_result[29]), .D(EX_ALU_result[28]), .Y(ALU__n123) );
  INVx1_ASAP7_75t_R ALU___U1767 ( .A(ALU__n1126), .Y(ALU__n1410) );
  NOR2x1p5_ASAP7_75t_R ALU___U1768 ( .A(EX_ALU_result[27]), .B(EX_ALU_result[26]), .Y(
        n1413) );
  NOR2x1p5_ASAP7_75t_R ALU___U1769 ( .A(EX_ALU_result[25]), .B(EX_ALU_result[24]), .Y(
        n1414) );
  INVx4_ASAP7_75t_R ALU___U1770 ( .A(ALU__n362), .Y(ALU__n1441) );
  INVx4_ASAP7_75t_R ALU___U1771 ( .A(ALU__n361), .Y(ALU__n1440) );
  BUFx12f_ASAP7_75t_R ALU___U1772 ( .A(ALU__n375), .Y(ALU__n1447) );
  BUFx5_ASAP7_75t_R ALU___U1773 ( .A(n1015), .Y(ALU__n1762) );
  BUFx5_ASAP7_75t_R ALU___U1774 ( .A(n1068), .Y(ALU__n1763) );
  BUFx5_ASAP7_75t_R ALU___U1775 ( .A(n1100), .Y(ALU__n1769) );
  BUFx5_ASAP7_75t_R ALU___U1776 ( .A(n920), .Y(ALU__n1771) );
  BUFx5_ASAP7_75t_R ALU___U1777 ( .A(n1060), .Y(ALU__n1776) );
  INVx5_ASAP7_75t_R ALU___U1778 ( .A(ALU__n1552), .Y(ALU__n1525) );
  BUFx6f_ASAP7_75t_R ALU___U1779 ( .A(ALU__n356), .Y(ALU__n1617) );
  BUFx12f_ASAP7_75t_R ALU___U1780 ( .A(ALU__n1426), .Y(ALU__n1616) );
  BUFx12f_ASAP7_75t_R ALU___U1781 ( .A(ALU__n1616), .Y(ALU__n1615) );
  BUFx3_ASAP7_75t_R ALU___U1782 ( .A(ALU__n1431), .Y(ALU__n1430) );
  BUFx2_ASAP7_75t_R ALU___U1783 ( .A(ALU__n329), .Y(ALU__n1431) );
  BUFx12f_ASAP7_75t_R ALU___U1784 ( .A(ALU__n986), .Y(ALU__n1644) );
  AND5x1_ASAP7_75t_R ALU___U1785 ( .A(ALU__n1620), .B(ALU__n1569), .C(ALU__n1309), .D(ALU__n1444), .E(
        n1506), .Y(ALU__n329) );
  BUFx16f_ASAP7_75t_R ALU___U1786 ( .A(ALU__n1193), .Y(ALU__n1569) );
  TIEHIx1_ASAP7_75t_R ALU___U1787 ( .H(ALU__n_Logic1_) );
  TIELOx1_ASAP7_75t_R ALU___U1788 ( .L(ALU__n6) );
  CKINVDCx14_ASAP7_75t_R ALU___U1789 ( .A(ALU__n844), .Y(ALU__n1432) );
  BUFx12f_ASAP7_75t_R ALU___U1790 ( .A(ALU__n1466), .Y(ALU__n1454) );
  BUFx12f_ASAP7_75t_R ALU___U1791 ( .A(ALU__n1163), .Y(ALU__n1459) );
  BUFx12f_ASAP7_75t_R ALU___U1792 ( .A(ALU__n1322), .Y(ALU__n1460) );
  BUFx12f_ASAP7_75t_R ALU___U1793 ( .A(ALU__n750), .Y(ALU__n1461) );
  BUFx12f_ASAP7_75t_R ALU___U1794 ( .A(ALU__n1321), .Y(ALU__n1462) );
  BUFx12f_ASAP7_75t_R ALU___U1795 ( .A(ALU__n1460), .Y(ALU__n1463) );
  CKINVDCx14_ASAP7_75t_R ALU___U1796 ( .A(ALU__n1507), .Y(ALU__n1505) );
  CKINVDCx14_ASAP7_75t_R ALU___U1797 ( .A(ALU__n1544), .Y(ALU__n1532) );
  CKINVDCx14_ASAP7_75t_R ALU___U1798 ( .A(ALU__n1541), .Y(ALU__n1535) );
  CKINVDCx14_ASAP7_75t_R ALU___U1799 ( .A(ALU__n1547), .Y(ALU__n1536) );
  CKINVDCx14_ASAP7_75t_R ALU___U1800 ( .A(ALU__n116), .Y(ALU__n1588) );
  OR2x2_ASAP7_75t_R ALU___U1801 ( .A(ALU__n1700), .B(n964), .Y(ALU__n1647) );
  OA21x2_ASAP7_75t_R ALU___U1802 ( .A1(ALU__n1053), .A2(n1015), .B(ALU__n1288), .Y(
        n1646) );
  OA221x2_ASAP7_75t_R ALU___U1803 ( .A1(ALU__n1746), .A2(n1060), .B1(ALU__n1683), 
        .B2(ALU__n1030), .C(ALU__n739), .Y(ALU__n1649) );
  OA221x2_ASAP7_75t_R ALU___U1804 ( .A1(ALU__n1682), .A2(n1233), .B1(ALU__n1747), 
        .B2(n1174), .C(ALU__n386), .Y(ALU__n1651) );
  OA221x2_ASAP7_75t_R ALU___U1805 ( .A1(ALU__n1235), .A2(n1114), .B1(ALU__n1194), 
        .B2(n973), .C(ALU__n388), .Y(ALU__n1653) );
  OA221x2_ASAP7_75t_R ALU___U1806 ( .A1(ALU__n903), .A2(n1029), .B1(ALU__n1680), 
        .B2(n929), .C(ALU__n407), .Y(ALU__n1655) );
  OA221x2_ASAP7_75t_R ALU___U1807 ( .A1(ALU__n1297), .A2(n1152), .B1(ALU__n1005), 
        .B2(n1229), .C(ALU__n673), .Y(ALU__n1657) );
  OA221x2_ASAP7_75t_R ALU___U1808 ( .A1(ALU__n1738), .A2(n1020), .B1(ALU__n1345), 
        .B2(n1109), .C(ALU__n670), .Y(ALU__n1659) );
  OA221x2_ASAP7_75t_R ALU___U1809 ( .A1(ALU__n1216), .A2(n925), .B1(ALU__n1697), 
        .B2(n969), .C(ALU__n848), .Y(ALU__n1661) );
  OA221x2_ASAP7_75t_R ALU___U1810 ( .A1(ALU__n1694), .A2(ALU__n965), .B1(ALU__n1695), .B2(
        n1073), .C(ALU__n766), .Y(ALU__n1663) );
  OA221x2_ASAP7_75t_R ALU___U1811 ( .A1(ALU__n1298), .A2(ALU__n904), .B1(ALU__n1065), .B2(
        n1182), .C(ALU__n768), .Y(ALU__n1665) );
  OA221x2_ASAP7_75t_R ALU___U1812 ( .A1(ALU__n1741), .A2(n1225), .B1(ALU__n1690), 
        .B2(n1068), .C(ALU__n427), .Y(ALU__n1667) );
  OA221x2_ASAP7_75t_R ALU___U1813 ( .A1(ALU__n1689), .A2(n1178), .B1(ALU__n1106), 
        .B2(n1024), .C(ALU__n735), .Y(ALU__n1669) );
  OA221x2_ASAP7_75t_R ALU___U1814 ( .A1(ALU__n1687), .A2(ALU__n934), .B1(ALU__n1688), .B2(
        n1064), .C(ALU__n733), .Y(ALU__n1671) );
  OA221x2_ASAP7_75t_R ALU___U1815 ( .A1(ALU__n1685), .A2(n1160), .B1(ALU__n1066), 
        .B2(n1100), .C(ALU__n621), .Y(ALU__n1673) );
  OA221x2_ASAP7_75t_R ALU___U1816 ( .A1(ALU__n938), .A2(n1215), .B1(ALU__n1105), 
        .B2(n920), .C(ALU__n892), .Y(ALU__n1675) );
  OA22x2_ASAP7_75t_R ALU___U1817 ( .A1(ALU__n691), .A2(ALU__n585), .B1(n888), .B2(
        n717), .Y(ALU__n1678) );
  INVx1_ASAP7_75t_R ALU___U1818 ( .A(n1222), .Y(ALU__n1740) );
  INVx1_ASAP7_75t_R ALU___U1819 ( .A(n619), .Y(ALU__n1749) );

  OAI311xp33_ASAP7_75t_R alu_control___U18 ( .A1(alu_control__alu_control__n167), .A2(inst_30_), .A3(alu_control__alu_control__n166), .B1(alu_control__n106), 
        .C1(alu_control__n48), .Y(alu_control__n16) );
  OA211x2_ASAP7_75t_R alu_control___U20 ( .A1(alu_control__n147), .A2(alu_control__n126), .B(alu_control__n135), .C(alu_control__n171), .Y(alu_control__n21)
         );
  OA22x2_ASAP7_75t_R alu_control___U21 ( .A1(alu_control__n147), .A2(alu_control__n116), .B1(alu_control__n173), .B2(alu_control__n85), .Y(alu_control__n20)
         );
  A2O1A1O1Ixp25_ASAP7_75t_R alu_control___U26 ( .A1(alu_control__n95), .A2(alu_control__n142), .B(alu_control__n133), .C(alu_control__n160), .D(
        n151), .Y(alu_control__n25) );
  OAI321xp33_ASAP7_75t_R alu_control___U28 ( .A1(alu_control__n155), .A2(alu_control__n120), .A3(alu_control__n154), .B1(alu_control__n167), 
        .B2(alu_control__n171), .C(alu_control__n156), .Y(alu_control__N106) );
  OR2x2_ASAP7_75t_R alu_control___U33 ( .A(inst_26_), .B(inst_25_), .Y(alu_control__n32) );
  OR2x2_ASAP7_75t_R alu_control___U37 ( .A(alu_control__n166), .B(alu_control__n65), .Y(alu_control__n18) );
  OR4x1_ASAP7_75t_R alu_control___U43 ( .A(inst_28_), .B(inst_27_), .C(inst_31_), .D(
        inst_29_), .Y(alu_control__n30) );
  DHLx3_ASAP7_75t_R alu_control___ALU_ctl_reg_3_ ( .CLK(alu_control__n152), .D(alu_control__n127), .Q(alu_control__n175) );
  DHLx3_ASAP7_75t_R alu_control___ALU_ctl_reg_2_ ( .CLK(alu_control__n152), .D(alu_control__n149), .Q(alu_control__n176) );
  DHLx3_ASAP7_75t_R alu_control___ALU_ctl_reg_1_ ( .CLK(alu_control__n152), .D(alu_control__n64), .Q(alu_control__n177) );
  DHLx3_ASAP7_75t_R alu_control___ALU_ctl_reg_0_ ( .CLK(alu_control__n152), .D(alu_control__n134), .Q(alu_control__n178) );
  HB1xp67_ASAP7_75t_R alu_control___U3 ( .A(alu_control__alu_control__n16), .Y(alu_control__n1) );
  HB1xp67_ASAP7_75t_R alu_control___U4 ( .A(alu_control__N106), .Y(alu_control__n2) );
  HB1xp67_ASAP7_75t_R alu_control___U5 ( .A(alu_control__n2), .Y(alu_control__n3) );
  HB1xp67_ASAP7_75t_R alu_control___U6 ( .A(alu_control__n3), .Y(alu_control__n4) );
  INVx13_ASAP7_75t_R alu_control___U7 ( .A(alu_control__n5), .Y(ALU_ctl[3]) );
  BUFx16f_ASAP7_75t_R alu_control___U8 ( .A(alu_control__n6), .Y(alu_control__n5) );
  BUFx12f_ASAP7_75t_R alu_control___U9 ( .A(alu_control__n102), .Y(alu_control__n6) );
  INVx5_ASAP7_75t_R alu_control___U10 ( .A(alu_control__n162), .Y(alu_control__n102) );
  BUFx4f_ASAP7_75t_R alu_control___U11 ( .A(alu_control__n28), .Y(alu_control__n7) );
  BUFx4f_ASAP7_75t_R alu_control___U12 ( .A(alu_control__n158), .Y(alu_control__n8) );
  BUFx3_ASAP7_75t_R alu_control___U13 ( .A(alu_control__n10), .Y(alu_control__n9) );
  BUFx2_ASAP7_75t_R alu_control___U14 ( .A(alu_control__n19), .Y(alu_control__n10) );
  BUFx2_ASAP7_75t_R alu_control___U15 ( .A(alu_control__n29), .Y(alu_control__n11) );
  AND3x1_ASAP7_75t_R alu_control___U16 ( .A(alu_control__n78), .B(alu_control__n57), .C(inst_13_), .Y(alu_control__n29) );
  BUFx12f_ASAP7_75t_R alu_control___U17 ( .A(alu_control__n176), .Y(alu_control__n12) );
  BUFx12f_ASAP7_75t_R alu_control___U19 ( .A(alu_control__n14), .Y(alu_control__n37) );
  INVx6_ASAP7_75t_R alu_control___U22 ( .A(alu_control__n55), .Y(alu_control__n159) );
  BUFx2_ASAP7_75t_R alu_control___U23 ( .A(alu_control__n41), .Y(alu_control__n38) );
  BUFx4f_ASAP7_75t_R alu_control___U24 ( .A(alu_control__n40), .Y(alu_control__n39) );
  BUFx3_ASAP7_75t_R alu_control___U25 ( .A(alu_control__n11), .Y(alu_control__n40) );
  BUFx2_ASAP7_75t_R alu_control___U27 ( .A(alu_control__n22), .Y(alu_control__n54) );
  INVx1_ASAP7_75t_R alu_control___U29 ( .A(alu_control__n54), .Y(alu_control__n41) );
  BUFx2_ASAP7_75t_R alu_control___U30 ( .A(alu_control__n71), .Y(alu_control__n42) );
  OR2x2_ASAP7_75t_R alu_control___U31 ( .A(alu_control__n69), .B(alu_control__n70), .Y(alu_control__n71) );
  BUFx2_ASAP7_75t_R alu_control___U32 ( .A(alu_control__n44), .Y(alu_control__n43) );
  BUFx2_ASAP7_75t_R alu_control___U34 ( .A(alu_control__n31), .Y(alu_control__n44) );
  BUFx2_ASAP7_75t_R alu_control___U35 ( .A(alu_control__n46), .Y(alu_control__n45) );
  BUFx2_ASAP7_75t_R alu_control___U36 ( .A(alu_control__n35), .Y(alu_control__n46) );
  BUFx2_ASAP7_75t_R alu_control___U38 ( .A(alu_control__n121), .Y(alu_control__n47) );
  AO22x2_ASAP7_75t_R alu_control___U39 ( .A1(alu_control__n157), .A2(alu_control__n58), .B1(alu_control__n160), .B2(alu_control__n47), .Y(alu_control__n31)
         );
  INVx1_ASAP7_75t_R alu_control___U40 ( .A(alu_control__n45), .Y(alu_control__n121) );
  BUFx6f_ASAP7_75t_R alu_control___U41 ( .A(alu_control__n49), .Y(alu_control__n48) );
  BUFx4f_ASAP7_75t_R alu_control___U42 ( .A(alu_control__n9), .Y(alu_control__n49) );
  OR2x2_ASAP7_75t_R alu_control___U44 ( .A(alu_control__n65), .B(alu_control__n79), .Y(alu_control__n19) );
  BUFx3_ASAP7_75t_R alu_control___U45 ( .A(alu_control__n51), .Y(alu_control__n50) );
  BUFx2_ASAP7_75t_R alu_control___U46 ( .A(alu_control__N108), .Y(alu_control__n51) );
  AO21x1_ASAP7_75t_R alu_control___U47 ( .A1(alu_control__n62), .A2(alu_control__n63), .B(alu_control__n159), .Y(alu_control__N108) );
  CKINVDCx16_ASAP7_75t_R alu_control___U48 ( .A(alu_control__n59), .Y(ALU_ctl[1]) );
  BUFx3_ASAP7_75t_R alu_control___U49 ( .A(alu_control__n53), .Y(alu_control__n52) );
  BUFx2_ASAP7_75t_R alu_control___U50 ( .A(alu_control__n36), .Y(alu_control__n53) );
  OR3x1_ASAP7_75t_R alu_control___U51 ( .A(inst_30_), .B(inst_13_), .C(alu_control__n142), .Y(alu_control__n36) );
  OR2x2_ASAP7_75t_R alu_control___U52 ( .A(alu_control__n68), .B(alu_control__n42), .Y(alu_control__n22) );
  BUFx12f_ASAP7_75t_R alu_control___U53 ( .A(alu_control__n56), .Y(alu_control__n55) );
  BUFx12f_ASAP7_75t_R alu_control___U54 ( .A(alu_control__n37), .Y(alu_control__n56) );
  BUFx3_ASAP7_75t_R alu_control___U55 ( .A(alu_control__n165), .Y(alu_control__n57) );
  BUFx2_ASAP7_75t_R alu_control___U56 ( .A(alu_control__n165), .Y(alu_control__n58) );
  INVx2_ASAP7_75t_R alu_control___U57 ( .A(inst_30_), .Y(alu_control__n165) );
  BUFx16f_ASAP7_75t_R alu_control___U58 ( .A(alu_control__n72), .Y(alu_control__n59) );
  BUFx12f_ASAP7_75t_R alu_control___U59 ( .A(alu_control__n83), .Y(alu_control__n72) );
  BUFx12f_ASAP7_75t_R alu_control___U60 ( .A(alu_control__n61), .Y(alu_control__n60) );
  BUFx12f_ASAP7_75t_R alu_control___U61 ( .A(alu_control__n17), .Y(alu_control__n61) );
  AO22x2_ASAP7_75t_R alu_control___U62 ( .A1(alu_control__n160), .A2(alu_control__n148), .B1(alu_control__n151), .B2(alu_control__n78), .Y(alu_control__n13)
         );
  INVx6_ASAP7_75t_R alu_control___U63 ( .A(alu_control__n60), .Y(alu_control__n151) );
  BUFx2_ASAP7_75t_R alu_control___U64 ( .A(alu_control__n20), .Y(alu_control__n62) );
  BUFx2_ASAP7_75t_R alu_control___U65 ( .A(alu_control__n21), .Y(alu_control__n63) );
  INVx1_ASAP7_75t_R alu_control___U66 ( .A(alu_control__n50), .Y(alu_control__n64) );
  BUFx3_ASAP7_75t_R alu_control___U67 ( .A(alu_control__n86), .Y(alu_control__n85) );
  BUFx6f_ASAP7_75t_R alu_control___U68 ( .A(alu_control__n66), .Y(alu_control__n65) );
  BUFx4f_ASAP7_75t_R alu_control___U69 ( .A(alu_control__n52), .Y(alu_control__n66) );
  BUFx3_ASAP7_75t_R alu_control___U70 ( .A(alu_control__n38), .Y(alu_control__n67) );
  INVx2_ASAP7_75t_R alu_control___U71 ( .A(inst_3_), .Y(alu_control__n69) );
  INVx3_ASAP7_75t_R alu_control___U72 ( .A(inst_2_), .Y(alu_control__n70) );
  INVx2_ASAP7_75t_R alu_control___U73 ( .A(alu_control__n136), .Y(alu_control__n68) );
  BUFx4f_ASAP7_75t_R alu_control___U74 ( .A(alu_control__n75), .Y(alu_control__n136) );
  BUFx3_ASAP7_75t_R alu_control___U75 ( .A(alu_control__n137), .Y(alu_control__n75) );
  INVx5_ASAP7_75t_R alu_control___U76 ( .A(alu_control__n145), .Y(alu_control__n83) );
  BUFx12f_ASAP7_75t_R alu_control___U77 ( .A(inst_14_), .Y(alu_control__n78) );
  BUFx6f_ASAP7_75t_R alu_control___U78 ( .A(alu_control__n74), .Y(alu_control__n73) );
  BUFx4f_ASAP7_75t_R alu_control___U79 ( .A(alu_control__n67), .Y(alu_control__n74) );
  BUFx12f_ASAP7_75t_R alu_control___U80 ( .A(alu_control__n178), .Y(alu_control__n76) );
  BUFx12f_ASAP7_75t_R alu_control___U81 ( .A(alu_control__n78), .Y(alu_control__n77) );
  BUFx6f_ASAP7_75t_R alu_control___U82 ( .A(inst_14_), .Y(alu_control__n79) );
  BUFx2_ASAP7_75t_R alu_control___U83 ( .A(alu_control__n26), .Y(alu_control__n80) );
  AND3x1_ASAP7_75t_R alu_control___U84 ( .A(alu_control__n115), .B(alu_control__n174), .C(inst_6_), .Y(alu_control__n26) );
  BUFx12f_ASAP7_75t_R alu_control___U85 ( .A(alu_control__n34), .Y(alu_control__n81) );
  INVx6_ASAP7_75t_R alu_control___U86 ( .A(alu_control__n140), .Y(alu_control__n157) );
  BUFx12f_ASAP7_75t_R alu_control___U87 ( .A(alu_control__n177), .Y(alu_control__n82) );
  INVx4_ASAP7_75t_R alu_control___U88 ( .A(alu_control__n77), .Y(alu_control__n166) );
  BUFx2_ASAP7_75t_R alu_control___U89 ( .A(alu_control__n23), .Y(alu_control__n86) );
  BUFx3_ASAP7_75t_R alu_control___U90 ( .A(alu_control__n88), .Y(alu_control__n87) );
  BUFx2_ASAP7_75t_R alu_control___U91 ( .A(alu_control__n24), .Y(alu_control__n88) );
  OR3x1_ASAP7_75t_R alu_control___U92 ( .A(inst_3_), .B(inst_6_), .C(inst_2_), .Y(alu_control__n24) );
  BUFx12f_ASAP7_75t_R alu_control___U93 ( .A(alu_control__N110), .Y(alu_control__n89) );
  AND2x4_ASAP7_75t_R alu_control___U94 ( .A(inst_30_), .B(alu_control__n8), .Y(alu_control__n28) );
  INVx2_ASAP7_75t_R alu_control___U95 ( .A(alu_control__n7), .Y(alu_control__n90) );
  AND2x4_ASAP7_75t_R alu_control___U96 ( .A(alu_control__n157), .B(alu_control__n166), .Y(alu_control__n158) );
  BUFx3_ASAP7_75t_R alu_control___U97 ( .A(alu_control__n92), .Y(alu_control__n91) );
  BUFx2_ASAP7_75t_R alu_control___U98 ( .A(alu_control__n18), .Y(alu_control__n92) );
  BUFx4f_ASAP7_75t_R alu_control___U99 ( .A(alu_control__n94), .Y(alu_control__n93) );
  BUFx3_ASAP7_75t_R alu_control___U100 ( .A(alu_control__n80), .Y(alu_control__n94) );
  INVx2_ASAP7_75t_R alu_control___U101 ( .A(alu_control__n125), .Y(alu_control__n174) );
  BUFx2_ASAP7_75t_R alu_control___U102 ( .A(alu_control__n96), .Y(alu_control__n95) );
  OA21x2_ASAP7_75t_R alu_control___U103 ( .A1(alu_control__n79), .A2(alu_control__n167), .B(alu_control__n106), .Y(alu_control__n23) );
  BUFx2_ASAP7_75t_R alu_control___U104 ( .A(alu_control__n143), .Y(alu_control__n164) );
  INVx1_ASAP7_75t_R alu_control___U105 ( .A(alu_control__n164), .Y(alu_control__n96) );
  BUFx3_ASAP7_75t_R alu_control___U106 ( .A(alu_control__n98), .Y(alu_control__n97) );
  BUFx2_ASAP7_75t_R alu_control___U107 ( .A(alu_control__n27), .Y(alu_control__n98) );
  BUFx3_ASAP7_75t_R alu_control___U108 ( .A(alu_control__n100), .Y(alu_control__n99) );
  BUFx2_ASAP7_75t_R alu_control___U109 ( .A(alu_control__N107), .Y(alu_control__n100) );
  INVx2_ASAP7_75t_R alu_control___U110 ( .A(alu_control__n39), .Y(alu_control__n143) );
  BUFx3_ASAP7_75t_R alu_control___U111 ( .A(alu_control__n132), .Y(alu_control__n131) );
  BUFx12f_ASAP7_75t_R alu_control___U112 ( .A(alu_control__n175), .Y(alu_control__n101) );
  BUFx6f_ASAP7_75t_R alu_control___U113 ( .A(alu_control__n105), .Y(alu_control__n104) );
  BUFx4f_ASAP7_75t_R alu_control___U114 ( .A(alu_control__n87), .Y(alu_control__n105) );
  BUFx6f_ASAP7_75t_R alu_control___U115 ( .A(alu_control__n107), .Y(alu_control__n106) );
  BUFx4f_ASAP7_75t_R alu_control___U116 ( .A(alu_control__n91), .Y(alu_control__n107) );
  BUFx2_ASAP7_75t_R alu_control___U117 ( .A(alu_control__n118), .Y(alu_control__n108) );
  BUFx2_ASAP7_75t_R alu_control___U118 ( .A(alu_control__n1), .Y(alu_control__alu_control__n109) );
  BUFx3_ASAP7_75t_R alu_control___U119 ( .A(alu_control__n111), .Y(alu_control__n110) );
  BUFx2_ASAP7_75t_R alu_control___U120 ( .A(alu_control__N109), .Y(alu_control__n111) );
  BUFx3_ASAP7_75t_R alu_control___U121 ( .A(alu_control__n113), .Y(alu_control__n112) );
  BUFx2_ASAP7_75t_R alu_control___U122 ( .A(alu_control__n13), .Y(alu_control__n113) );
  BUFx4f_ASAP7_75t_R alu_control___U123 ( .A(inst_5_), .Y(alu_control__n114) );
  BUFx2_ASAP7_75t_R alu_control___U124 ( .A(inst_5_), .Y(alu_control__n115) );
  BUFx2_ASAP7_75t_R alu_control___U125 ( .A(inst_5_), .Y(alu_control__n116) );
  BUFx3_ASAP7_75t_R alu_control___U126 ( .A(alu_control__n108), .Y(alu_control__n117) );
  BUFx2_ASAP7_75t_R alu_control___U127 ( .A(alu_control__n4), .Y(alu_control__n118) );
  BUFx2_ASAP7_75t_R alu_control___U128 ( .A(alu_control__n33), .Y(alu_control__n119) );
  AO21x1_ASAP7_75t_R alu_control___U129 ( .A1(alu_control__n171), .A2(alu_control__n173), .B(alu_control__n159), .Y(alu_control__n33) );
  INVx1_ASAP7_75t_R alu_control___U130 ( .A(alu_control__n43), .Y(alu_control__n120) );
  AND4x1_ASAP7_75t_R alu_control___U131 ( .A(alu_control__n90), .B(alu_control__n106), .C(alu_control__n48), .D(alu_control__n143), .Y(alu_control__n35) );
  BUFx6f_ASAP7_75t_R alu_control___U132 ( .A(inst_12_), .Y(alu_control__n122) );
  BUFx4f_ASAP7_75t_R alu_control___U133 ( .A(inst_12_), .Y(alu_control__n123) );
  BUFx3_ASAP7_75t_R alu_control___U134 ( .A(inst_4_), .Y(alu_control__n124) );
  BUFx4f_ASAP7_75t_R alu_control___U135 ( .A(inst_4_), .Y(alu_control__n125) );
  BUFx2_ASAP7_75t_R alu_control___U136 ( .A(inst_4_), .Y(alu_control__n126) );
  OR2x6_ASAP7_75t_R alu_control___U137 ( .A(alu_control__n159), .B(alu_control__n135), .Y(alu_control__N110) );
  INVx6_ASAP7_75t_R alu_control___U138 ( .A(alu_control__n89), .Y(alu_control__n127) );
  INVx2_ASAP7_75t_R alu_control___U139 ( .A(alu_control__n127), .Y(alu_control__n169) );
  INVx3_ASAP7_75t_R alu_control___U140 ( .A(alu_control__n104), .Y(alu_control__n128) );
  AND3x4_ASAP7_75t_R alu_control___U141 ( .A(alu_control__n128), .B(alu_control__n114), .C(alu_control__n124), .Y(alu_control__n15) );
  BUFx4f_ASAP7_75t_R alu_control___U142 ( .A(alu_control__n128), .Y(alu_control__n172) );
  BUFx12f_ASAP7_75t_R alu_control___U143 ( .A(alu_control__n130), .Y(ALU_ctl[0]) );
  BUFx12f_ASAP7_75t_R alu_control___U144 ( .A(alu_control__n76), .Y(alu_control__n130) );
  BUFx2_ASAP7_75t_R alu_control___U145 ( .A(alu_control__n25), .Y(alu_control__n132) );
  AND2x2_ASAP7_75t_R alu_control___U146 ( .A(alu_control__n90), .B(alu_control__n48), .Y(alu_control__n27) );
  INVx1_ASAP7_75t_R alu_control___U147 ( .A(alu_control__n97), .Y(alu_control__n133) );
  OA21x2_ASAP7_75t_R alu_control___U148 ( .A1(alu_control__n131), .A2(alu_control__n159), .B(alu_control__n169), .Y(alu_control__N107) );
  INVx1_ASAP7_75t_R alu_control___U149 ( .A(alu_control__n99), .Y(alu_control__n134) );
  INVx3_ASAP7_75t_R alu_control___U150 ( .A(alu_control__n73), .Y(alu_control__n135) );
  BUFx2_ASAP7_75t_R alu_control___U151 ( .A(alu_control__n144), .Y(alu_control__n170) );
  INVx1_ASAP7_75t_R alu_control___U152 ( .A(alu_control__n170), .Y(alu_control__n137) );
  BUFx12f_ASAP7_75t_R alu_control___U153 ( .A(alu_control__n139), .Y(ALU_ctl[2]) );
  BUFx12f_ASAP7_75t_R alu_control___U154 ( .A(alu_control__n12), .Y(alu_control__n139) );
  BUFx12f_ASAP7_75t_R alu_control___U155 ( .A(alu_control__n141), .Y(alu_control__n140) );
  BUFx12f_ASAP7_75t_R alu_control___U156 ( .A(alu_control__n81), .Y(alu_control__n141) );
  OR2x6_ASAP7_75t_R alu_control___U157 ( .A(alu_control__n123), .B(inst_13_), .Y(alu_control__n34) );
  BUFx6f_ASAP7_75t_R alu_control___U158 ( .A(alu_control__n122), .Y(alu_control__n168) );
  INVx3_ASAP7_75t_R alu_control___U159 ( .A(alu_control__n168), .Y(alu_control__n142) );
  INVx3_ASAP7_75t_R alu_control___U160 ( .A(alu_control__n151), .Y(alu_control__n171) );
  INVx2_ASAP7_75t_R alu_control___U161 ( .A(alu_control__n93), .Y(alu_control__n144) );
  BUFx16f_ASAP7_75t_R alu_control___U162 ( .A(alu_control__n146), .Y(alu_control__n145) );
  BUFx12f_ASAP7_75t_R alu_control___U163 ( .A(alu_control__n82), .Y(alu_control__n146) );
  INVx2_ASAP7_75t_R alu_control___U164 ( .A(alu_control__n172), .Y(alu_control__n147) );
  BUFx2_ASAP7_75t_R alu_control___U165 ( .A(alu_control__n109), .Y(alu_control__n148) );
  OA21x2_ASAP7_75t_R alu_control___U166 ( .A1(alu_control__n150), .A2(alu_control__n159), .B(alu_control__n169), .Y(alu_control__N109) );
  INVx1_ASAP7_75t_R alu_control___U167 ( .A(alu_control__n110), .Y(alu_control__n149) );
  INVx1_ASAP7_75t_R alu_control___U168 ( .A(alu_control__n112), .Y(alu_control__n150) );
  OR3x2_ASAP7_75t_R alu_control___U169 ( .A(inst_3_), .B(inst_2_), .C(alu_control__n144), .Y(alu_control__n17) );
  BUFx6f_ASAP7_75t_R alu_control___U170 ( .A(alu_control__n153), .Y(alu_control__n152) );
  BUFx4f_ASAP7_75t_R alu_control___U171 ( .A(alu_control__n117), .Y(alu_control__n153) );
  BUFx2_ASAP7_75t_R alu_control___U172 ( .A(alu_control__n32), .Y(alu_control__n154) );
  BUFx2_ASAP7_75t_R alu_control___U173 ( .A(alu_control__n30), .Y(alu_control__n155) );
  INVx1_ASAP7_75t_R alu_control___U174 ( .A(alu_control__n119), .Y(alu_control__n156) );
  INVx3_ASAP7_75t_R alu_control___U175 ( .A(alu_control__n157), .Y(alu_control__n167) );
  AND2x6_ASAP7_75t_R alu_control___U176 ( .A(inst_1_), .B(inst_0_), .Y(alu_control__n14) );
  BUFx12f_ASAP7_75t_R alu_control___U177 ( .A(alu_control__n161), .Y(alu_control__n160) );
  BUFx12f_ASAP7_75t_R alu_control___U178 ( .A(alu_control__n15), .Y(alu_control__n161) );
  INVx3_ASAP7_75t_R alu_control___U179 ( .A(alu_control__n160), .Y(alu_control__n173) );
  BUFx16f_ASAP7_75t_R alu_control___U180 ( .A(alu_control__n163), .Y(alu_control__n162) );
  BUFx12f_ASAP7_75t_R alu_control___U181 ( .A(alu_control__n101), .Y(alu_control__n163) );

 BUFx5_ASAP7_75t_R CONTROL_HAZARD_U1 ( .A(Branch), .Y(IF_flush) );
BUFx5_ASAP7_75t_R CONTROL_HAZARD_U2 ( .A(ALU_zero), .Y(ID_flush) );
 XOR2x2_ASAP7_75t_R EX_DW01_add_1___U2 ( .A(EX_DW01_add_1__n205), .B(EX_DW01_add_1__n232), .Y(EX_branch_addr[7]) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U3 ( .A(EX_DW01_add_1__n407), .B(EX_DW01_add_1__n544), .Y(EX_DW01_add_1__n540) );
  AND3x2_ASAP7_75t_R EX_DW01_add_1___U4 ( .A(EX_DW01_add_1__n47), .B(EX_DW01_add_1__n18), .C(EX_DW01_add_1__n616), .Y(EX_DW01_add_1__n153) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U5 ( .A(EX_DW01_add_1__EX_DW01_add_1__n153), .Y(EX_DW01_add_1__n1) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U6 ( .A(EX_DW01_add_1__n153), .Y(EX_DW01_add_1__n2) );
  BUFx16f_ASAP7_75t_R EX_DW01_add_1___U7 ( .A(EX_DW01_add_1__n404), .Y(EX_DW01_add_1__n3) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U8 ( .A(EX_DW01_add_1__n405), .Y(EX_DW01_add_1__n404) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U9 ( .A(EX_DW01_add_1__n190), .Y(EX_DW01_add_1__n57) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U10 ( .A(EX_DW01_add_1__n287), .Y(EX_DW01_add_1__n62) );
  NAND2x1p5_ASAP7_75t_R EX_DW01_add_1___U11 ( .A(ID_EX_imm[4]), .B(inst_addr[4]), .Y(EX_DW01_add_1__n40) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U12 ( .A(ID_EX_imm[23]), .B(inst_addr[23]), .Y(EX_DW01_add_1__n567) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U13 ( .A(EX_DW01_add_1__n361), .Y(EX_DW01_add_1__n469) );
  BUFx16f_ASAP7_75t_R EX_DW01_add_1___U14 ( .A(EX_DW01_add_1__n362), .Y(EX_DW01_add_1__n361) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U15 ( .A(EX_DW01_add_1__n226), .Y(EX_DW01_add_1__n370) );
  BUFx16f_ASAP7_75t_R EX_DW01_add_1___U16 ( .A(EX_DW01_add_1__n227), .Y(EX_DW01_add_1__n226) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U17 ( .A(EX_DW01_add_1__n224), .Y(EX_DW01_add_1__n366) );
  BUFx16f_ASAP7_75t_R EX_DW01_add_1___U18 ( .A(EX_DW01_add_1__n225), .Y(EX_DW01_add_1__n224) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U19 ( .A(EX_DW01_add_1__n229), .Y(EX_DW01_add_1__n351) );
  BUFx16f_ASAP7_75t_R EX_DW01_add_1___U20 ( .A(EX_DW01_add_1__n230), .Y(EX_DW01_add_1__n229) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U21 ( .A(EX_DW01_add_1__n174), .Y(EX_DW01_add_1__n207) );
  BUFx16f_ASAP7_75t_R EX_DW01_add_1___U22 ( .A(EX_DW01_add_1__n175), .Y(EX_DW01_add_1__n174) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U23 ( .A(EX_DW01_add_1__n106), .Y(EX_DW01_add_1__n393) );
  NOR2xp67_ASAP7_75t_R EX_DW01_add_1___U24 ( .A(EX_DW01_add_1__n116), .B(EX_DW01_add_1__n123), .Y(EX_DW01_add_1__n70) );
  NOR2x1_ASAP7_75t_R EX_DW01_add_1___U25 ( .A(inst_addr[15]), .B(ID_EX_imm[15]), .Y(EX_DW01_add_1__n123) );
  NAND2xp67_ASAP7_75t_R EX_DW01_add_1___U26 ( .A(ID_EX_imm[15]), .B(inst_addr[15]), .Y(EX_DW01_add_1__n67) );
  NAND2x1p5_ASAP7_75t_R EX_DW01_add_1___U27 ( .A(EX_DW01_add_1__n329), .B(EX_DW01_add_1__n568), .Y(EX_DW01_add_1__n117) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U28 ( .A(EX_DW01_add_1__n329), .B(EX_DW01_add_1__n568), .Y(EX_DW01_add_1__n13) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U29 ( .A(EX_DW01_add_1__n5), .Y(EX_DW01_add_1__n4) );
  AOI21xp33_ASAP7_75t_R EX_DW01_add_1___U30 ( .A1(EX_DW01_add_1__n151), .A2(EX_DW01_add_1__n68), .B(EX_DW01_add_1__n354), .Y(EX_DW01_add_1__n5) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U31 ( .A(EX_DW01_add_1__n139), .B(EX_DW01_add_1__n147), .Y(EX_branch_addr[6]) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U32 ( .A(ID_EX_imm[22]), .Y(EX_DW01_add_1__n6) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U33 ( .A(EX_DW01_add_1__n583), .B(EX_DW01_add_1__n217), .Y(EX_branch_addr[21]) );
  NOR2x1_ASAP7_75t_R EX_DW01_add_1___U34 ( .A(EX_DW01_add_1__n313), .B(EX_DW01_add_1__n464), .Y(EX_DW01_add_1__n7) );
  NOR2x1p5_ASAP7_75t_R EX_DW01_add_1___U35 ( .A(EX_DW01_add_1__n7), .B(EX_DW01_add_1__n477), .Y(EX_DW01_add_1__n411) );
  INVx4_ASAP7_75t_R EX_DW01_add_1___U36 ( .A(EX_DW01_add_1__n504), .Y(EX_DW01_add_1__n464) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U37 ( .A(EX_DW01_add_1__n668), .Y(EX_branch_addr[4]) );
  INVx6_ASAP7_75t_R EX_DW01_add_1___U38 ( .A(EX_DW01_add_1__n298), .Y(EX_DW01_add_1__n129) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U39 ( .A(EX_DW01_add_1__n5), .Y(EX_DW01_add_1__n8) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U40 ( .A(EX_DW01_add_1__n565), .Y(EX_DW01_add_1__n480) );
  INVx4_ASAP7_75t_R EX_DW01_add_1___U41 ( .A(EX_DW01_add_1__n336), .Y(EX_DW01_add_1__n447) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U42 ( .A(EX_DW01_add_1__n447), .Y(EX_DW01_add_1__n497) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U43 ( .A(EX_DW01_add_1__n432), .B(EX_DW01_add_1__n447), .Y(EX_DW01_add_1__n498) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U44 ( .A(EX_DW01_add_1__n644), .B(EX_DW01_add_1__n89), .Y(EX_DW01_add_1__n9) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U45 ( .A(EX_DW01_add_1__EX_DW01_add_1__n108), .Y(EX_DW01_add_1__n10) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U46 ( .A(EX_DW01_add_1__n9), .B(EX_DW01_add_1__n10), .Y(EX_DW01_add_1__EX_DW01_add_1__n109) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U47 ( .A(EX_DW01_add_1__n486), .B(EX_DW01_add_1__n379), .Y(EX_DW01_add_1__n89) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U48 ( .A(EX_DW01_add_1__n349), .B(EX_DW01_add_1__n429), .Y(EX_DW01_add_1__n108) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U49 ( .A(EX_DW01_add_1__n109), .B(EX_DW01_add_1__n66), .Y(EX_DW01_add_1__n61) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U50 ( .A(EX_DW01_add_1__n346), .Y(EX_DW01_add_1__n11) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U51 ( .A(EX_DW01_add_1__n140), .B(EX_DW01_add_1__n152), .Y(EX_DW01_add_1__n313) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U52 ( .A(EX_DW01_add_1__n329), .B(EX_DW01_add_1__n568), .Y(EX_DW01_add_1__n12) );
  AND3x1_ASAP7_75t_R EX_DW01_add_1___U53 ( .A(EX_DW01_add_1__n59), .B(EX_DW01_add_1__n371), .C(EX_DW01_add_1__n400), .Y(EX_DW01_add_1__n14) );
  AND3x1_ASAP7_75t_R EX_DW01_add_1___U54 ( .A(EX_DW01_add_1__n59), .B(EX_DW01_add_1__n371), .C(EX_DW01_add_1__n400), .Y(EX_DW01_add_1__n15) );
  A2O1A1Ixp33_ASAP7_75t_R EX_DW01_add_1___U55 ( .A1(EX_DW01_add_1__n28), .A2(EX_DW01_add_1__n450), .B(EX_DW01_add_1__n11), .C(EX_DW01_add_1__n368), .Y(EX_DW01_add_1__n16) );
  OAI21x1_ASAP7_75t_R EX_DW01_add_1___U56 ( .A1(EX_DW01_add_1__n316), .A2(EX_DW01_add_1__n375), .B(EX_DW01_add_1__EX_DW01_add_1__n281), .Y(EX_DW01_add_1__n28) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U57 ( .A(EX_DW01_add_1__n620), .Y(EX_DW01_add_1__n17) );
  NAND3xp33_ASAP7_75t_R EX_DW01_add_1___U58 ( .A(EX_DW01_add_1__n47), .B(EX_DW01_add_1__n18), .C(EX_DW01_add_1__n616), .Y(EX_DW01_add_1__n39) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U59 ( .A(EX_DW01_add_1__n15), .B(EX_DW01_add_1__n617), .Y(EX_DW01_add_1__n18) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U60 ( .A(EX_DW01_add_1__n46), .Y(EX_DW01_add_1__n617) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U61 ( .A(EX_DW01_add_1__n280), .B(EX_DW01_add_1__n655), .Y(EX_DW01_add_1__n79) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U62 ( .A(EX_DW01_add_1__n412), .B(EX_DW01_add_1__n432), .Y(EX_DW01_add_1__n655) );
  NAND2x1p5_ASAP7_75t_R EX_DW01_add_1___U63 ( .A(EX_DW01_add_1__n128), .B(EX_DW01_add_1__n408), .Y(EX_DW01_add_1__n152) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U64 ( .A(EX_DW01_add_1__n422), .Y(EX_DW01_add_1__n268) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U65 ( .A(EX_DW01_add_1__n533), .B(EX_DW01_add_1__n295), .Y(EX_DW01_add_1__n136) );
  NAND2x1p5_ASAP7_75t_R EX_DW01_add_1___U66 ( .A(EX_DW01_add_1__n647), .B(EX_DW01_add_1__n617), .Y(EX_DW01_add_1__n54) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U67 ( .A(EX_DW01_add_1__n432), .Y(EX_DW01_add_1__n431) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U68 ( .A(EX_DW01_add_1__n38), .Y(EX_DW01_add_1__n432) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U69 ( .A(EX_DW01_add_1__n19), .B(EX_DW01_add_1__n20), .Y(EX_branch_addr[15]) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U70 ( .A(EX_DW01_add_1__n207), .Y(EX_DW01_add_1__n19) );
  AOI21xp5_ASAP7_75t_R EX_DW01_add_1___U71 ( .A1(EX_DW01_add_1__n71), .A2(EX_DW01_add_1__n623), .B(EX_DW01_add_1__n471), .Y(EX_DW01_add_1__n20) );
  NAND2x1p5_ASAP7_75t_R EX_DW01_add_1___U72 ( .A(EX_DW01_add_1__n141), .B(EX_DW01_add_1__n49), .Y(EX_DW01_add_1__n94) );
  NAND2xp67_ASAP7_75t_R EX_DW01_add_1___U73 ( .A(EX_DW01_add_1__n283), .B(EX_DW01_add_1__n95), .Y(EX_DW01_add_1__n46) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U74 ( .A(EX_DW01_add_1__n94), .Y(EX_DW01_add_1__n95) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U75 ( .A(EX_DW01_add_1__n116), .Y(EX_DW01_add_1__n471) );
  NAND2x1p5_ASAP7_75t_R EX_DW01_add_1___U76 ( .A(ID_EX_imm[14]), .B(inst_addr[14]), .Y(EX_DW01_add_1__n116) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U77 ( .A(EX_DW01_add_1__n620), .Y(EX_DW01_add_1__n382) );
  NOR2x1p5_ASAP7_75t_R EX_DW01_add_1___U78 ( .A(EX_DW01_add_1__n80), .B(EX_DW01_add_1__n79), .Y(EX_DW01_add_1__n620) );
  NOR2x1_ASAP7_75t_R EX_DW01_add_1___U79 ( .A(EX_DW01_add_1__n122), .B(EX_DW01_add_1__n620), .Y(EX_DW01_add_1__n639) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U80 ( .A(EX_DW01_add_1__n119), .B(EX_DW01_add_1__n87), .Y(EX_DW01_add_1__n120) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U81 ( .A(EX_DW01_add_1__n15), .Y(EX_DW01_add_1__n21) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U82 ( .A(EX_DW01_add_1__n525), .Y(EX_DW01_add_1__n300) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U83 ( .A(EX_DW01_add_1__n300), .Y(EX_DW01_add_1__n299) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U84 ( .A(EX_DW01_add_1__n503), .Y(EX_DW01_add_1__n412) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U85 ( .A(EX_DW01_add_1__n61), .B(EX_DW01_add_1__n60), .Y(EX_DW01_add_1__n154) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U86 ( .A(EX_DW01_add_1__n66), .B(EX_DW01_add_1__n109), .Y(EX_DW01_add_1__n75) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U87 ( .A(EX_DW01_add_1__n487), .Y(EX_DW01_add_1__n308) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U88 ( .A(EX_DW01_add_1__n656), .Y(EX_DW01_add_1__n381) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U89 ( .A(inst_addr[7]), .B(ID_EX_imm[7]), .Y(EX_DW01_add_1__n496) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U90 ( .A(EX_DW01_add_1__n412), .Y(EX_DW01_add_1__n500) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U91 ( .A(EX_DW01_add_1__n540), .Y(EX_DW01_add_1__n426) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U92 ( .A(EX_DW01_add_1__n557), .Y(EX_DW01_add_1__n85) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U93 ( .A(EX_DW01_add_1__n330), .Y(EX_DW01_add_1__n329) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U94 ( .A(EX_DW01_add_1__n140), .B(EX_DW01_add_1__n152), .Y(EX_DW01_add_1__n22) );
  AOI21xp33_ASAP7_75t_R EX_DW01_add_1___U95 ( .A1(EX_DW01_add_1__n515), .A2(EX_DW01_add_1__n115), .B(EX_DW01_add_1__n97), .Y(EX_DW01_add_1__n517) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U96 ( .A(EX_DW01_add_1__n115), .B(EX_DW01_add_1__n34), .Y(EX_DW01_add_1__n103) );
  AOI21xp5_ASAP7_75t_R EX_DW01_add_1___U97 ( .A1(EX_DW01_add_1__n639), .A2(EX_DW01_add_1__n333), .B(EX_DW01_add_1__n289), .Y(EX_DW01_add_1__n133) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U98 ( .A(EX_DW01_add_1__n488), .Y(EX_DW01_add_1__n445) );
  NAND2x1p5_ASAP7_75t_R EX_DW01_add_1___U99 ( .A(ID_EX_imm[5]), .B(inst_addr[5]), .Y(EX_DW01_add_1__n42) );
  AND3x1_ASAP7_75t_R EX_DW01_add_1___U100 ( .A(EX_DW01_add_1__n462), .B(EX_DW01_add_1__n396), .C(EX_DW01_add_1__n653), .Y(EX_DW01_add_1__n408) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U101 ( .A(EX_DW01_add_1__n475), .Y(EX_DW01_add_1__n304) );
  AOI21x1_ASAP7_75t_R EX_DW01_add_1___U102 ( .A1(EX_DW01_add_1__n480), .A2(EX_DW01_add_1__n30), .B(EX_DW01_add_1__n144), .Y(EX_DW01_add_1__n24) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U103 ( .A(EX_DW01_add_1__n23), .B(EX_DW01_add_1__n228), .Y(EX_DW01_add_1__n663) );
  NAND2xp67_ASAP7_75t_R EX_DW01_add_1___U104 ( .A(EX_DW01_add_1__n377), .B(EX_DW01_add_1__n142), .Y(EX_DW01_add_1__n23) );
  INVx6_ASAP7_75t_R EX_DW01_add_1___U105 ( .A(EX_DW01_add_1__n299), .Y(EX_DW01_add_1__n467) );
  OAI21xp5_ASAP7_75t_R EX_DW01_add_1___U106 ( .A1(EX_DW01_add_1__n398), .A2(EX_DW01_add_1__n416), .B(EX_DW01_add_1__n298), .Y(EX_DW01_add_1__n81) );
  XNOR2xp5_ASAP7_75t_R EX_DW01_add_1___U107 ( .A(EX_DW01_add_1__n88), .B(EX_DW01_add_1__n24), .Y(EX_DW01_add_1__n659) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U108 ( .A(EX_DW01_add_1__n423), .Y(EX_DW01_add_1__n25) );
  NAND2x1_ASAP7_75t_R EX_DW01_add_1___U109 ( .A(EX_DW01_add_1__n451), .B(EX_DW01_add_1__n83), .Y(EX_DW01_add_1__n142) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U110 ( .A(EX_DW01_add_1__n353), .B(EX_DW01_add_1__n623), .Y(EX_DW01_add_1__n26) );
  NAND3xp33_ASAP7_75t_R EX_DW01_add_1___U111 ( .A(EX_DW01_add_1__n27), .B(EX_DW01_add_1__n49), .C(EX_DW01_add_1__n283), .Y(EX_DW01_add_1__n72) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U112 ( .A(EX_DW01_add_1__n26), .Y(EX_DW01_add_1__n27) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U113 ( .A(EX_DW01_add_1__n627), .Y(EX_DW01_add_1__n353) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U114 ( .A(EX_DW01_add_1__n120), .B(EX_DW01_add_1__n435), .Y(EX_DW01_add_1__n557) );
  NAND2x1_ASAP7_75t_R EX_DW01_add_1___U115 ( .A(EX_DW01_add_1__n43), .B(EX_DW01_add_1__n84), .Y(EX_DW01_add_1__n100) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U116 ( .A(ID_EX_imm[11]), .B(inst_addr[11]), .Y(EX_DW01_add_1__n645) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U117 ( .A(EX_DW01_add_1__n117), .Y(EX_DW01_add_1__n29) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U118 ( .A(EX_DW01_add_1__n568), .Y(EX_DW01_add_1__n30) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U119 ( .A(EX_DW01_add_1__n12), .Y(EX_DW01_add_1__n555) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U120 ( .A(EX_DW01_add_1__n320), .Y(EX_DW01_add_1__n319) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U121 ( .A(EX_DW01_add_1__n349), .B(EX_DW01_add_1__n429), .Y(EX_DW01_add_1__n32) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U122 ( .A(EX_DW01_add_1__n624), .Y(EX_DW01_add_1__n383) );
  NAND3xp33_ASAP7_75t_R EX_DW01_add_1___U123 ( .A(EX_DW01_add_1__EX_DW01_add_1__n154), .B(EX_DW01_add_1__n1), .C(EX_DW01_add_1__EX_DW01_add_1__n104), .Y(EX_DW01_add_1__n31) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U124 ( .A(EX_DW01_add_1__n574), .Y(EX_DW01_add_1__n375) );
  NAND2xp67_ASAP7_75t_R EX_DW01_add_1___U125 ( .A(EX_DW01_add_1__n377), .B(EX_DW01_add_1__n41), .Y(EX_DW01_add_1__n71) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U126 ( .A(EX_DW01_add_1__n640), .Y(EX_DW01_add_1__n413) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U127 ( .A(EX_DW01_add_1__n347), .Y(EX_DW01_add_1__n346) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U128 ( .A(EX_DW01_add_1__n252), .B(EX_DW01_add_1__n552), .Y(EX_DW01_add_1__n45) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U129 ( .A(EX_DW01_add_1__n515), .B(EX_DW01_add_1__n372), .Y(EX_DW01_add_1__n33) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U130 ( .A(EX_DW01_add_1__n33), .Y(EX_DW01_add_1__n34) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U131 ( .A(EX_DW01_add_1__n373), .Y(EX_DW01_add_1__n372) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U132 ( .A(inst_addr[22]), .Y(EX_DW01_add_1__n35) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U133 ( .A(EX_DW01_add_1__n178), .B(EX_DW01_add_1__n36), .Y(EX_branch_addr[17]) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U134 ( .A(EX_DW01_add_1__n96), .Y(EX_DW01_add_1__n36) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U135 ( .A(EX_DW01_add_1__n561), .Y(EX_DW01_add_1__n435) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U136 ( .A(EX_DW01_add_1__n192), .B(EX_DW01_add_1__n37), .Y(EX_branch_addr[18]) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U137 ( .A(EX_DW01_add_1__n98), .Y(EX_DW01_add_1__n37) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U138 ( .A(inst_addr[6]), .B(ID_EX_imm[6]), .Y(EX_DW01_add_1__n38) );
  NAND3xp33_ASAP7_75t_R EX_DW01_add_1___U139 ( .A(EX_DW01_add_1__n100), .B(EX_DW01_add_1__n135), .C(EX_DW01_add_1__n332), .Y(EX_DW01_add_1__n47) );
  NOR2x1_ASAP7_75t_R EX_DW01_add_1___U140 ( .A(EX_DW01_add_1__n51), .B(EX_DW01_add_1__n50), .Y(EX_DW01_add_1__n527) );
  NOR2x1_ASAP7_75t_R EX_DW01_add_1___U141 ( .A(EX_DW01_add_1__n53), .B(EX_DW01_add_1__n45), .Y(EX_DW01_add_1__n50) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U142 ( .A(EX_DW01_add_1__n348), .Y(EX_DW01_add_1__n118) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U143 ( .A(EX_DW01_add_1__n105), .B(EX_DW01_add_1__n609), .Y(EX_DW01_add_1__n422) );
  OAI21x1_ASAP7_75t_R EX_DW01_add_1___U144 ( .A1(EX_DW01_add_1__n473), .A2(EX_DW01_add_1__n411), .B(EX_DW01_add_1__n42), .Y(EX_DW01_add_1__n139) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U145 ( .A(EX_DW01_add_1__n136), .Y(EX_DW01_add_1__n521) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U146 ( .A(EX_DW01_add_1__n451), .B(EX_DW01_add_1__n83), .Y(EX_DW01_add_1__n41) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U147 ( .A(EX_DW01_add_1__n82), .Y(EX_DW01_add_1__n83) );
  XOR2x2_ASAP7_75t_R EX_DW01_add_1___U148 ( .A(EX_DW01_add_1__n206), .B(EX_DW01_add_1__n485), .Y(EX_branch_addr[9]) );
  NAND2xp67_ASAP7_75t_R EX_DW01_add_1___U149 ( .A(EX_DW01_add_1__n374), .B(EX_DW01_add_1__n103), .Y(EX_DW01_add_1__n63) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U150 ( .A(EX_DW01_add_1__n353), .B(EX_DW01_add_1__n623), .Y(EX_DW01_add_1__n141) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U151 ( .A(EX_DW01_add_1__n279), .B(EX_DW01_add_1__n129), .Y(EX_DW01_add_1__n43) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U152 ( .A(EX_DW01_add_1__n128), .B(EX_DW01_add_1__n408), .Y(EX_DW01_add_1__n44) );
  NAND2x1p5_ASAP7_75t_R EX_DW01_add_1___U153 ( .A(EX_DW01_add_1__n283), .B(EX_DW01_add_1__n95), .Y(EX_DW01_add_1__n438) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U154 ( .A(EX_DW01_add_1__n481), .Y(EX_DW01_add_1__n618) );
  INVx4_ASAP7_75t_R EX_DW01_add_1___U155 ( .A(EX_DW01_add_1__n319), .Y(EX_DW01_add_1__n481) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U156 ( .A(EX_DW01_add_1__n481), .Y(EX_DW01_add_1__n616) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U157 ( .A(EX_DW01_add_1__n116), .B(EX_DW01_add_1__n123), .Y(EX_DW01_add_1__n48) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U158 ( .A(EX_DW01_add_1__n471), .Y(EX_DW01_add_1__n322) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U159 ( .A(inst_addr[15]), .B(ID_EX_imm[15]), .Y(EX_DW01_add_1__n49) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U160 ( .A(EX_DW01_add_1__n235), .Y(EX_DW01_add_1__n51) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U161 ( .A(EX_DW01_add_1__n67), .Y(EX_DW01_add_1__n441) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U162 ( .A(EX_DW01_add_1__n67), .Y(EX_DW01_add_1__n479) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U163 ( .A(EX_DW01_add_1__n252), .B(EX_DW01_add_1__n552), .Y(EX_DW01_add_1__n115) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U164 ( .A(EX_DW01_add_1__n127), .B(EX_DW01_add_1__n56), .Y(EX_branch_addr[27]) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U165 ( .A(inst_addr[28]), .B(ID_EX_imm[28]), .Y(EX_DW01_add_1__n534) );
  NAND3x1_ASAP7_75t_R EX_DW01_add_1___U166 ( .A(EX_DW01_add_1__n2), .B(EX_DW01_add_1__n154), .C(EX_DW01_add_1__n104), .Y(EX_DW01_add_1__n52) );
  NAND3x1_ASAP7_75t_R EX_DW01_add_1___U167 ( .A(EX_DW01_add_1__n154), .B(EX_DW01_add_1__n39), .C(EX_DW01_add_1__n104), .Y(EX_DW01_add_1__n151) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U168 ( .A(EX_DW01_add_1__n438), .Y(EX_DW01_add_1__n619) );
  OAI21xp5_ASAP7_75t_R EX_DW01_add_1___U169 ( .A1(EX_DW01_add_1__n548), .A2(EX_DW01_add_1__n45), .B(EX_DW01_add_1__n326), .Y(EX_DW01_add_1__n64) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U170 ( .A(EX_DW01_add_1__n521), .Y(EX_DW01_add_1__n53) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U171 ( .A(EX_DW01_add_1__n595), .Y(EX_DW01_add_1__n279) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U172 ( .A(EX_DW01_add_1__n14), .B(EX_DW01_add_1__n22), .Y(EX_DW01_add_1__n640) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U173 ( .A(EX_DW01_add_1__n517), .B(EX_DW01_add_1__n55), .Y(EX_branch_addr[30]) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U174 ( .A(EX_DW01_add_1__n114), .Y(EX_DW01_add_1__n55) );
  NOR2x2_ASAP7_75t_R EX_DW01_add_1___U175 ( .A(EX_DW01_add_1__n542), .B(EX_DW01_add_1__n326), .Y(EX_DW01_add_1__n92) );
  OAI21xp5_ASAP7_75t_R EX_DW01_add_1___U176 ( .A1(EX_DW01_add_1__n304), .A2(EX_DW01_add_1__n45), .B(EX_DW01_add_1__n417), .Y(EX_DW01_add_1__n107) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U177 ( .A(EX_DW01_add_1__n476), .B(EX_DW01_add_1__n273), .Y(EX_DW01_add_1__n533) );
  INVx4_ASAP7_75t_R EX_DW01_add_1___U178 ( .A(EX_DW01_add_1__n277), .Y(EX_DW01_add_1__n326) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U179 ( .A(EX_DW01_add_1__n632), .Y(EX_DW01_add_1__n451) );
  OAI21xp5_ASAP7_75t_R EX_DW01_add_1___U180 ( .A1(EX_DW01_add_1__n426), .A2(EX_DW01_add_1__n45), .B(EX_DW01_add_1__n355), .Y(EX_DW01_add_1__n56) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U181 ( .A(inst_addr[13]), .B(ID_EX_imm[13]), .Y(EX_DW01_add_1__n627) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U182 ( .A(ID_EX_imm[13]), .B(inst_addr[13]), .Y(EX_DW01_add_1__n402) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U183 ( .A(EX_DW01_add_1__n57), .B(EX_DW01_add_1__n527), .Y(EX_branch_addr[29]) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U184 ( .A(EX_DW01_add_1__n75), .B(EX_DW01_add_1__n121), .Y(EX_DW01_add_1__n110) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U185 ( .A(ID_EX_imm[6]), .B(inst_addr[6]), .Y(EX_DW01_add_1__n499) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U186 ( .A(EX_DW01_add_1__n432), .B(EX_DW01_add_1__n412), .Y(EX_DW01_add_1__n59) );
  OA21x2_ASAP7_75t_R EX_DW01_add_1___U187 ( .A1(EX_DW01_add_1__n398), .A2(EX_DW01_add_1__n416), .B(EX_DW01_add_1__n298), .Y(EX_DW01_add_1__n58) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U188 ( .A(EX_DW01_add_1__n467), .Y(EX_DW01_add_1__n298) );
  INVx3_ASAP7_75t_R EX_DW01_add_1___U189 ( .A(EX_DW01_add_1__n524), .Y(EX_DW01_add_1__n416) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U190 ( .A(EX_DW01_add_1__n65), .Y(EX_DW01_add_1__n66) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U191 ( .A(EX_DW01_add_1__n44), .B(EX_DW01_add_1__n113), .Y(EX_DW01_add_1__n125) );
  AND3x4_ASAP7_75t_R EX_DW01_add_1___U192 ( .A(EX_DW01_add_1__n59), .B(EX_DW01_add_1__n371), .C(EX_DW01_add_1__n400), .Y(EX_DW01_add_1__n647) );
  NAND3xp33_ASAP7_75t_R EX_DW01_add_1___U193 ( .A(EX_DW01_add_1__n17), .B(EX_DW01_add_1__n91), .C(EX_DW01_add_1__n618), .Y(EX_DW01_add_1__n60) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U194 ( .A(EX_DW01_add_1__n90), .Y(EX_DW01_add_1__n91) );
  AOI21xp5_ASAP7_75t_R EX_DW01_add_1___U195 ( .A1(EX_DW01_add_1__n644), .A2(EX_DW01_add_1__n89), .B(EX_DW01_add_1__n32), .Y(EX_DW01_add_1__n624) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U196 ( .A(inst_addr[0]), .B(n731), .Y(EX_DW01_add_1__n595) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U197 ( .A(EX_DW01_add_1__n62), .B(EX_DW01_add_1__n63), .Y(EX_branch_addr[31]) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U198 ( .A(EX_DW01_add_1__n295), .Y(EX_DW01_add_1__n529) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U199 ( .A(EX_DW01_add_1__n532), .Y(EX_DW01_add_1__n294) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U200 ( .A(EX_DW01_add_1__n394), .Y(EX_DW01_add_1__n274) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U201 ( .A(EX_DW01_add_1__n619), .B(EX_DW01_add_1__n625), .Y(EX_DW01_add_1__n65) );
  AOI22xp5_ASAP7_75t_R EX_DW01_add_1___U202 ( .A1(EX_DW01_add_1__n553), .A2(EX_DW01_add_1__n329), .B1(EX_DW01_add_1__n29), .B2(EX_DW01_add_1__n137), .Y(
        n126) );
  NOR2x1p5_ASAP7_75t_R EX_DW01_add_1___U203 ( .A(EX_DW01_add_1__n590), .B(EX_DW01_add_1__n143), .Y(EX_DW01_add_1__n137) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U204 ( .A(EX_DW01_add_1__n42), .Y(EX_DW01_add_1__n502) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U205 ( .A(EX_DW01_add_1__n588), .Y(EX_DW01_add_1__n354) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U206 ( .A(EX_DW01_add_1__n267), .B(EX_DW01_add_1__n334), .Y(EX_DW01_add_1__n68) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U207 ( .A(inst_addr[16]), .Y(EX_DW01_add_1__n69) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U208 ( .A(EX_DW01_add_1__n267), .B(EX_DW01_add_1__n334), .Y(EX_DW01_add_1__n558) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U209 ( .A(EX_DW01_add_1__n249), .Y(EX_DW01_add_1__n119) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U210 ( .A(EX_DW01_add_1__n133), .B(EX_DW01_add_1__n111), .Y(EX_DW01_add_1__n485) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U211 ( .A(EX_DW01_add_1__n654), .Y(EX_DW01_add_1__n280) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U212 ( .A(EX_DW01_add_1__n619), .B(EX_DW01_add_1__n400), .Y(EX_DW01_add_1__n90) );
  NOR2x1p5_ASAP7_75t_R EX_DW01_add_1___U213 ( .A(EX_DW01_add_1__n77), .B(EX_DW01_add_1__n325), .Y(EX_DW01_add_1__n73) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U214 ( .A(EX_DW01_add_1__n78), .Y(EX_DW01_add_1__n74) );
  NOR2x2_ASAP7_75t_R EX_DW01_add_1___U215 ( .A(EX_DW01_add_1__n74), .B(EX_DW01_add_1__n73), .Y(EX_DW01_add_1__n590) );
  INVx4_ASAP7_75t_R EX_DW01_add_1___U216 ( .A(EX_DW01_add_1__n599), .Y(EX_DW01_add_1__n77) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U217 ( .A(EX_DW01_add_1__n265), .Y(EX_DW01_add_1__n78) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U218 ( .A(ID_EX_imm[24]), .B(inst_addr[24]), .Y(EX_DW01_add_1__n563) );
  NOR3x1_ASAP7_75t_R EX_DW01_add_1___U219 ( .A(EX_DW01_add_1__n638), .B(EX_DW01_add_1__n425), .C(EX_DW01_add_1__n640), .Y(EX_DW01_add_1__n632) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U220 ( .A(EX_DW01_add_1__n5), .Y(EX_DW01_add_1__n76) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U221 ( .A(EX_DW01_add_1__n343), .B(EX_DW01_add_1__n353), .Y(EX_DW01_add_1__n82) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U222 ( .A(EX_DW01_add_1__n325), .Y(EX_DW01_add_1__n478) );
  NOR2x1_ASAP7_75t_R EX_DW01_add_1___U223 ( .A(EX_DW01_add_1__n143), .B(EX_DW01_add_1__n590), .Y(EX_DW01_add_1__n315) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U224 ( .A(EX_DW01_add_1__n381), .Y(EX_DW01_add_1__n80) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U225 ( .A(EX_DW01_add_1__n601), .Y(EX_DW01_add_1__n325) );
  OAI21x1_ASAP7_75t_R EX_DW01_add_1___U226 ( .A1(EX_DW01_add_1__n485), .A2(EX_DW01_add_1__n397), .B(EX_DW01_add_1__n307), .Y(EX_DW01_add_1__n146) );
  NAND2x1p5_ASAP7_75t_R EX_DW01_add_1___U227 ( .A(EX_DW01_add_1__n350), .B(EX_DW01_add_1__n396), .Y(EX_DW01_add_1__n135) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U228 ( .A(EX_DW01_add_1__n332), .B(EX_DW01_add_1__n396), .Y(EX_DW01_add_1__n507) );
  AND3x1_ASAP7_75t_R EX_DW01_add_1___U229 ( .A(EX_DW01_add_1__n462), .B(EX_DW01_add_1__n396), .C(EX_DW01_add_1__n653), .Y(EX_DW01_add_1__n84) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U230 ( .A(EX_DW01_add_1__n638), .Y(EX_DW01_add_1__n436) );
  OAI21xp5_ASAP7_75t_R EX_DW01_add_1___U231 ( .A1(EX_DW01_add_1__n485), .A2(EX_DW01_add_1__n397), .B(EX_DW01_add_1__n307), .Y(EX_DW01_add_1__n99) );
  AOI21xp5_ASAP7_75t_R EX_DW01_add_1___U232 ( .A1(EX_DW01_add_1__n99), .A2(EX_DW01_add_1__n379), .B(EX_DW01_add_1__n474), .Y(EX_DW01_add_1__n132) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U233 ( .A(EX_DW01_add_1__n409), .Y(EX_DW01_add_1__n88) );
  O2A1O1Ixp5_ASAP7_75t_R EX_DW01_add_1___U234 ( .A1(EX_DW01_add_1__n535), .A2(EX_DW01_add_1__n92), .B(EX_DW01_add_1__n274), .C(EX_DW01_add_1__n537), .Y(
        n130) );
  OAI21xp5_ASAP7_75t_R EX_DW01_add_1___U235 ( .A1(EX_DW01_add_1__n519), .A2(EX_DW01_add_1__n101), .B(EX_DW01_add_1__n102), .Y(EX_DW01_add_1__n516) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U236 ( .A(EX_DW01_add_1__n346), .B(EX_DW01_add_1__n423), .Y(EX_DW01_add_1__n568) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U237 ( .A(EX_DW01_add_1__n72), .B(EX_DW01_add_1__n118), .Y(EX_DW01_add_1__n86) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U238 ( .A(EX_DW01_add_1__n86), .Y(EX_DW01_add_1__n87) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U239 ( .A(EX_DW01_add_1__n590), .Y(EX_DW01_add_1__n428) );
  AND3x1_ASAP7_75t_R EX_DW01_add_1___U240 ( .A(EX_DW01_add_1__n89), .B(EX_DW01_add_1__n625), .C(EX_DW01_add_1__n333), .Y(EX_DW01_add_1__n320) );
  NAND3xp33_ASAP7_75t_R EX_DW01_add_1___U241 ( .A(EX_DW01_add_1__n91), .B(EX_DW01_add_1__n382), .C(EX_DW01_add_1__n618), .Y(EX_DW01_add_1__n121) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U242 ( .A(EX_DW01_add_1__n646), .Y(EX_DW01_add_1__n379) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U243 ( .A(EX_DW01_add_1__n555), .Y(EX_DW01_add_1__n93) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U244 ( .A(EX_DW01_add_1__n602), .Y(EX_DW01_add_1__n599) );
  O2A1O1Ixp33_ASAP7_75t_R EX_DW01_add_1___U245 ( .A1(EX_DW01_add_1__n535), .A2(EX_DW01_add_1__n92), .B(EX_DW01_add_1__n273), .C(EX_DW01_add_1__n537), .Y(
        n530) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U246 ( .A(EX_DW01_add_1__n461), .B(EX_DW01_add_1__n281), .Y(EX_DW01_add_1__n423) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U247 ( .A(EX_DW01_add_1__n366), .Y(EX_DW01_add_1__n96) );
  OAI21xp33_ASAP7_75t_R EX_DW01_add_1___U248 ( .A1(EX_DW01_add_1__n519), .A2(EX_DW01_add_1__n101), .B(EX_DW01_add_1__n102), .Y(EX_DW01_add_1__n97) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U249 ( .A(EX_DW01_add_1__n390), .Y(EX_DW01_add_1__n101) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U250 ( .A(ID_EX_imm[9]), .B(inst_addr[9]), .Y(EX_DW01_add_1__n487) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U251 ( .A(EX_DW01_add_1__n469), .Y(EX_DW01_add_1__n98) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U252 ( .A(EX_DW01_add_1__n251), .Y(EX_DW01_add_1__n284) );
  OAI31xp33_ASAP7_75t_R EX_DW01_add_1___U253 ( .A1(EX_DW01_add_1__n85), .A2(EX_DW01_add_1__n556), .A3(EX_DW01_add_1__n110), .B(EX_DW01_add_1__n558), .Y(
        n150) );
  NAND2xp67_ASAP7_75t_R EX_DW01_add_1___U254 ( .A(ID_EX_imm[29]), .B(inst_addr[29]), .Y(EX_DW01_add_1__n102) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U255 ( .A(EX_DW01_add_1__n394), .Y(EX_DW01_add_1__n273) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U256 ( .A(EX_DW01_add_1__n395), .Y(EX_DW01_add_1__n394) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U257 ( .A(EX_DW01_add_1__n652), .Y(EX_DW01_add_1__n111) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U258 ( .A(EX_DW01_add_1__n449), .Y(EX_DW01_add_1__n537) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U259 ( .A(EX_DW01_add_1__n271), .Y(EX_DW01_add_1__n395) );
  INVxp67_ASAP7_75t_R EX_DW01_add_1___U260 ( .A(EX_DW01_add_1__n302), .Y(EX_DW01_add_1__n374) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U261 ( .A(EX_DW01_add_1__n513), .Y(EX_DW01_add_1__n302) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U262 ( .A(EX_DW01_add_1__n272), .Y(EX_DW01_add_1__n271) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U263 ( .A(EX_DW01_add_1__n621), .B(EX_DW01_add_1__n561), .Y(EX_DW01_add_1__n104) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U264 ( .A(EX_DW01_add_1__n536), .Y(EX_DW01_add_1__n272) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U265 ( .A(EX_DW01_add_1__n519), .Y(EX_DW01_add_1__n235) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U266 ( .A(EX_DW01_add_1__n602), .B(EX_DW01_add_1__n610), .Y(EX_DW01_add_1__n105) );
  NAND2xp5_ASAP7_75t_R EX_DW01_add_1___U267 ( .A(EX_DW01_add_1__n609), .B(EX_DW01_add_1__n610), .Y(EX_DW01_add_1__n106) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U268 ( .A(EX_DW01_add_1__n599), .Y(EX_DW01_add_1__n352) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U269 ( .A(EX_DW01_add_1__n265), .Y(EX_DW01_add_1__n399) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U270 ( .A(EX_DW01_add_1__n199), .B(EX_DW01_add_1__n107), .Y(EX_branch_addr[28]) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U271 ( .A(EX_DW01_add_1__n58), .B(EX_DW01_add_1__n233), .Y(EX_DW01_add_1__n670) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U272 ( .A(EX_DW01_add_1__n509), .Y(EX_DW01_add_1__n276) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U273 ( .A(EX_DW01_add_1__n670), .Y(EX_branch_addr[2]) );
  INVx4_ASAP7_75t_R EX_DW01_add_1___U274 ( .A(EX_DW01_add_1__n453), .Y(EX_DW01_add_1__n526) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U275 ( .A(EX_DW01_add_1__n413), .Y(EX_DW01_add_1__n259) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U276 ( .A(EX_DW01_add_1__n194), .B(EX_DW01_add_1__n508), .Y(EX_DW01_add_1__n669) );
  NAND2xp33_ASAP7_75t_R EX_DW01_add_1___U277 ( .A(EX_DW01_add_1__n135), .B(EX_DW01_add_1__n332), .Y(EX_DW01_add_1__n112) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U278 ( .A(EX_DW01_add_1__n112), .Y(EX_DW01_add_1__n113) );
  INVx4_ASAP7_75t_R EX_DW01_add_1___U279 ( .A(EX_DW01_add_1__n337), .Y(EX_DW01_add_1__n446) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U280 ( .A(EX_DW01_add_1__n446), .Y(EX_DW01_add_1__n339) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U281 ( .A(EX_DW01_add_1__n138), .Y(EX_DW01_add_1__n114) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U282 ( .A(EX_DW01_add_1__n468), .Y(EX_DW01_add_1__n492) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U283 ( .A(EX_DW01_add_1__n666), .Y(EX_branch_addr[8]) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U284 ( .A(EX_DW01_add_1__n669), .Y(EX_branch_addr[3]) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U285 ( .A(EX_DW01_add_1__n49), .Y(EX_DW01_add_1__n629) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U286 ( .A(n762), .B(inst_addr[3]), .Y(EX_DW01_add_1__n510) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U287 ( .A(EX_DW01_add_1__n635), .B(EX_DW01_add_1__n444), .Y(EX_branch_addr[13]) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U288 ( .A(EX_DW01_add_1__n641), .B(EX_DW01_add_1__n406), .Y(EX_DW01_add_1__n664) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U289 ( .A(EX_DW01_add_1__n135), .B(EX_DW01_add_1__n332), .Y(EX_DW01_add_1__n140) );
  AOI21x1_ASAP7_75t_R EX_DW01_add_1___U290 ( .A1(EX_DW01_add_1__n456), .A2(EX_DW01_add_1__n189), .B(EX_DW01_add_1__n269), .Y(EX_DW01_add_1__n601) );
  INVx3_ASAP7_75t_R EX_DW01_add_1___U291 ( .A(EX_DW01_add_1__n456), .Y(EX_DW01_add_1__n472) );
  CKINVDCx5p33_ASAP7_75t_R EX_DW01_add_1___U292 ( .A(EX_DW01_add_1__n189), .Y(EX_DW01_add_1__n455) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U293 ( .A(EX_DW01_add_1__n269), .Y(EX_DW01_add_1__n414) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U294 ( .A(EX_DW01_add_1__n664), .Y(EX_branch_addr[12]) );
  XNOR2xp5_ASAP7_75t_R EX_DW01_add_1___U295 ( .A(EX_DW01_add_1__n445), .B(EX_DW01_add_1__n392), .Y(EX_DW01_add_1__n666) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U296 ( .A(EX_DW01_add_1__n639), .Y(EX_DW01_add_1__n468) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U297 ( .A(EX_DW01_add_1__n146), .B(EX_DW01_add_1__n218), .Y(EX_DW01_add_1__n665) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U298 ( .A(EX_DW01_add_1__n306), .Y(EX_DW01_add_1__n410) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U299 ( .A(EX_DW01_add_1__n306), .Y(EX_DW01_add_1__n305) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U300 ( .A(EX_DW01_add_1__n661), .Y(EX_branch_addr[19]) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U301 ( .A(EX_DW01_add_1__n586), .Y(EX_DW01_add_1__n306) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U302 ( .A(EX_DW01_add_1__n446), .Y(EX_DW01_add_1__n349) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U303 ( .A(EX_DW01_add_1__n663), .Y(EX_branch_addr[14]) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U304 ( .A(EX_DW01_add_1__n400), .Y(EX_DW01_add_1__n122) );
  AOI21x1_ASAP7_75t_R EX_DW01_add_1___U305 ( .A1(EX_DW01_add_1__n68), .A2(EX_DW01_add_1__n151), .B(EX_DW01_add_1__n354), .Y(EX_DW01_add_1__n565) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U306 ( .A(EX_DW01_add_1__n4), .B(EX_DW01_add_1__n124), .Y(EX_DW01_add_1__n660) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U307 ( .A(EX_DW01_add_1__n351), .Y(EX_DW01_add_1__n124) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U308 ( .A(EX_DW01_add_1__n660), .Y(EX_branch_addr[20]) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U309 ( .A(EX_DW01_add_1__n449), .B(EX_DW01_add_1__n273), .Y(EX_DW01_add_1__n127) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U310 ( .A(EX_DW01_add_1__n349), .Y(EX_DW01_add_1__n474) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U311 ( .A(EX_DW01_add_1__n279), .B(EX_DW01_add_1__n129), .Y(EX_DW01_add_1__n128) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U312 ( .A(EX_DW01_add_1__n284), .Y(EX_DW01_add_1__n283) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U313 ( .A(EX_DW01_add_1__n418), .Y(EX_DW01_add_1__n417) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U314 ( .A(EX_DW01_add_1__n345), .B(EX_DW01_add_1__n64), .Y(EX_branch_addr[26]) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U315 ( .A(EX_DW01_add_1__n131), .B(EX_DW01_add_1__n132), .Y(EX_branch_addr[11]) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U316 ( .A(EX_DW01_add_1__n134), .Y(EX_DW01_add_1__n131) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U317 ( .A(EX_DW01_add_1__n492), .Y(EX_DW01_add_1__n425) );
  XNOR2xp5_ASAP7_75t_R EX_DW01_add_1___U318 ( .A(EX_DW01_add_1__EX_DW01_add_1__n459), .B(EX_DW01_add_1__n45), .Y(EX_branch_addr[25]) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U319 ( .A(EX_DW01_add_1__n667), .Y(EX_branch_addr[5]) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U320 ( .A(EX_DW01_add_1__n370), .Y(EX_DW01_add_1__n134) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U321 ( .A(EX_DW01_add_1__n357), .Y(EX_DW01_add_1__n439) );
  INVxp33_ASAP7_75t_R EX_DW01_add_1___U322 ( .A(EX_DW01_add_1__n439), .Y(EX_DW01_add_1__n475) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U323 ( .A(ID_EX_imm[2]), .B(inst_addr[2]), .Y(EX_DW01_add_1__n523) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U324 ( .A(EX_DW01_add_1__n596), .Y(EX_DW01_add_1__n181) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U325 ( .A(EX_DW01_add_1__n181), .B(EX_DW01_add_1__n231), .Y(EX_DW01_add_1__n661) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U326 ( .A(EX_DW01_add_1__n16), .Y(EX_DW01_add_1__n144) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U327 ( .A(EX_DW01_add_1__n559), .Y(EX_DW01_add_1__n348) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U328 ( .A(EX_DW01_add_1__n452), .Y(EX_DW01_add_1__n290) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U329 ( .A(ID_EX_imm[8]), .B(inst_addr[8]), .Y(EX_DW01_add_1__n452) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U330 ( .A(EX_DW01_add_1__n348), .Y(EX_DW01_add_1__n483) );
  AND3x1_ASAP7_75t_R EX_DW01_add_1___U331 ( .A(EX_DW01_add_1__n623), .B(EX_DW01_add_1__n49), .C(EX_DW01_add_1__n402), .Y(EX_DW01_add_1__n559) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U332 ( .A(EX_DW01_add_1__n560), .Y(EX_DW01_add_1__n246) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U333 ( .A(EX_DW01_add_1__n625), .B(EX_DW01_add_1__n383), .Y(EX_DW01_add_1__n638) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U334 ( .A(EX_DW01_add_1__n246), .Y(EX_DW01_add_1__n250) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U335 ( .A(EX_DW01_add_1__n250), .Y(EX_DW01_add_1__n249) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U336 ( .A(ID_EX_imm[26]), .B(inst_addr[26]), .Y(EX_DW01_add_1__n545) );
  AO22x1_ASAP7_75t_R EX_DW01_add_1___U337 ( .A1(ID_EX_imm[30]), .A2(inst_addr[30]), .B1(EX_DW01_add_1__n372), .B2(EX_DW01_add_1__n516), .Y(
        n513) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U338 ( .A(EX_DW01_add_1__n3), .Y(EX_DW01_add_1__n138) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U339 ( .A(EX_DW01_add_1__n344), .Y(EX_DW01_add_1__n418) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U340 ( .A(EX_DW01_add_1__n544), .Y(EX_DW01_add_1__n542) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U341 ( .A(EX_DW01_add_1__n530), .Y(EX_DW01_add_1__n344) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U342 ( .A(ID_EX_imm[12]), .B(inst_addr[12]), .Y(EX_DW01_add_1__n622) );
  XNOR2xp5_ASAP7_75t_R EX_DW01_add_1___U343 ( .A(EX_DW01_add_1__n411), .B(EX_DW01_add_1__n424), .Y(EX_DW01_add_1__n667) );
  XNOR2xp5_ASAP7_75t_R EX_DW01_add_1___U344 ( .A(EX_DW01_add_1__n313), .B(EX_DW01_add_1__n442), .Y(EX_DW01_add_1__n668) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U345 ( .A(inst_addr[1]), .B(ID_EX_imm[1]), .Y(EX_DW01_add_1__n525) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U346 ( .A(inst_addr[11]), .B(ID_EX_imm[11]), .Y(EX_DW01_add_1__n625) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U347 ( .A(EX_DW01_add_1__n546), .Y(EX_DW01_add_1__n407) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U348 ( .A(EX_DW01_add_1__n581), .Y(EX_DW01_add_1__n340) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U349 ( .A(EX_DW01_add_1__n544), .B(EX_DW01_add_1__n430), .Y(EX_DW01_add_1__n547) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U350 ( .A(EX_DW01_add_1__n539), .Y(EX_DW01_add_1__n476) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U351 ( .A(EX_DW01_add_1__n623), .B(EX_DW01_add_1__n322), .Y(EX_DW01_add_1__n630) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U352 ( .A(EX_DW01_add_1__n426), .Y(EX_DW01_add_1__n539) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U353 ( .A(EX_DW01_add_1__n440), .Y(EX_DW01_add_1__n357) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U354 ( .A(EX_DW01_add_1__n358), .Y(EX_DW01_add_1__n440) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U355 ( .A(EX_DW01_add_1__n533), .Y(EX_DW01_add_1__n358) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U356 ( .A(ID_EX_imm[8]), .B(inst_addr[8]), .Y(EX_DW01_add_1__n491) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U357 ( .A(EX_DW01_add_1__n491), .Y(EX_DW01_add_1__n333) );
  CKINVDCx20_ASAP7_75t_R EX_DW01_add_1___U358 ( .A(EX_DW01_add_1__n334), .Y(EX_DW01_add_1__n143) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U359 ( .A(EX_DW01_add_1__n610), .Y(EX_DW01_add_1__n606) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U360 ( .A(ID_EX_imm[26]), .B(inst_addr[26]), .Y(EX_DW01_add_1__n544) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U361 ( .A(EX_DW01_add_1__n234), .Y(EX_DW01_add_1__n145) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U362 ( .A(EX_DW01_add_1__n145), .Y(EX_DW01_add_1__n147) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U363 ( .A(EX_DW01_add_1__n6), .B(EX_DW01_add_1__n35), .Y(EX_DW01_add_1__n566) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U364 ( .A(ID_EX_imm[5]), .B(inst_addr[5]), .Y(EX_DW01_add_1__n503) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U365 ( .A(n2), .B(ID_EX_imm[21]), .Y(EX_DW01_add_1__n581) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U366 ( .A(inst_addr[9]), .B(ID_EX_imm[9]), .Y(EX_DW01_add_1__n486) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U367 ( .A(inst_addr[14]), .B(ID_EX_imm[14]), .Y(EX_DW01_add_1__n623) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U368 ( .A(n1), .B(ID_EX_imm[25]), .Y(EX_DW01_add_1__n546) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U369 ( .A(EX_DW01_add_1__n461), .Y(EX_DW01_add_1__n285) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U370 ( .A(EX_DW01_add_1__n582), .B(EX_DW01_add_1__n340), .Y(EX_DW01_add_1__n461) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U371 ( .A(EX_DW01_add_1__n493), .Y(EX_DW01_add_1__n205) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U372 ( .A(EX_DW01_add_1__n275), .Y(EX_DW01_add_1__n463) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U373 ( .A(ID_EX_imm[7]), .B(inst_addr[7]), .Y(EX_DW01_add_1__n427) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U374 ( .A(EX_DW01_add_1__n576), .B(EX_DW01_add_1__n367), .Y(EX_branch_addr[22]) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U375 ( .A(ID_EX_imm[17]), .B(inst_addr[17]), .Y(EX_DW01_add_1__n608) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U376 ( .A(ID_EX_imm[20]), .Y(EX_DW01_add_1__n148) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U377 ( .A(inst_addr[20]), .Y(EX_DW01_add_1__n149) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U378 ( .A(EX_DW01_add_1__n148), .B(EX_DW01_add_1__n149), .Y(EX_DW01_add_1__n586) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U379 ( .A(EX_DW01_add_1__n665), .Y(EX_branch_addr[10]) );
  XOR2xp5_ASAP7_75t_R EX_DW01_add_1___U380 ( .A(EX_DW01_add_1__n443), .B(EX_DW01_add_1__n570), .Y(EX_branch_addr[23]) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U381 ( .A(EX_DW01_add_1__n453), .Y(EX_DW01_add_1__n657) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U382 ( .A(EX_DW01_add_1__n279), .Y(EX_DW01_add_1__n342) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U383 ( .A(EX_DW01_add_1__n499), .Y(EX_DW01_add_1__n336) );
  INVx6_ASAP7_75t_R EX_DW01_add_1___U384 ( .A(EX_DW01_add_1__n341), .Y(EX_DW01_add_1__n453) );
  HB1xp67_ASAP7_75t_R EX_DW01_add_1___U385 ( .A(EX_DW01_add_1__n659), .Y(EX_branch_addr[24]) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U386 ( .A(inst_addr[10]), .B(ID_EX_imm[10]), .Y(EX_DW01_add_1__n646) );
  XNOR2xp5_ASAP7_75t_R EX_DW01_add_1___U387 ( .A(EX_DW01_add_1__n369), .B(EX_DW01_add_1__n52), .Y(EX_DW01_add_1__n662) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U388 ( .A(EX_DW01_add_1__n628), .Y(EX_DW01_add_1__n155) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U389 ( .A(EX_DW01_add_1__n501), .Y(EX_DW01_add_1__n156) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U390 ( .A(EX_DW01_add_1__n494), .Y(EX_DW01_add_1__n157) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U391 ( .A(EX_DW01_add_1__n400), .Y(EX_DW01_add_1__n495) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U392 ( .A(EX_DW01_add_1__n577), .Y(EX_DW01_add_1__n158) );
  AO21x1_ASAP7_75t_R EX_DW01_add_1___U393 ( .A1(EX_DW01_add_1__n582), .A2(EX_DW01_add_1__n8), .B(EX_DW01_add_1__n410), .Y(EX_DW01_add_1__n583) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U394 ( .A(EX_DW01_add_1__n160), .Y(EX_DW01_add_1__n159) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U395 ( .A(EX_DW01_add_1__n672), .Y(EX_DW01_add_1__n160) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U396 ( .A(EX_DW01_add_1__n484), .Y(EX_DW01_add_1__n161) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U397 ( .A(EX_DW01_add_1__n522), .Y(EX_DW01_add_1__n162) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U398 ( .A(EX_DW01_add_1__n611), .Y(EX_DW01_add_1__n163) );
  AO21x1_ASAP7_75t_R EX_DW01_add_1___U399 ( .A1(EX_DW01_add_1__n31), .A2(EX_DW01_add_1__n609), .B(EX_DW01_add_1__n614), .Y(EX_DW01_add_1__n611) );
  AO21x1_ASAP7_75t_R EX_DW01_add_1___U400 ( .A1(EX_DW01_add_1__n480), .A2(EX_DW01_add_1__n285), .B(EX_DW01_add_1__n193), .Y(EX_DW01_add_1__n576) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U401 ( .A(EX_DW01_add_1__n165), .Y(EX_DW01_add_1__n164) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U402 ( .A(EX_DW01_add_1__n156), .Y(EX_DW01_add_1__n165) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U403 ( .A(EX_DW01_add_1__n502), .B(EX_DW01_add_1__n473), .Y(EX_DW01_add_1__n501) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U404 ( .A(EX_DW01_add_1__n615), .Y(EX_DW01_add_1__n166) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U405 ( .A(EX_DW01_add_1__n612), .Y(EX_DW01_add_1__n167) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U406 ( .A(EX_DW01_add_1__n603), .Y(EX_DW01_add_1__n168) );
  AO21x1_ASAP7_75t_R EX_DW01_add_1___U407 ( .A1(EX_DW01_add_1__n52), .A2(EX_DW01_add_1__n393), .B(EX_DW01_add_1__n478), .Y(EX_DW01_add_1__n603) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U408 ( .A(EX_DW01_add_1__n648), .Y(EX_DW01_add_1__n169) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U409 ( .A(EX_DW01_add_1__n636), .Y(EX_DW01_add_1__n170) );
  AND3x1_ASAP7_75t_R EX_DW01_add_1___U410 ( .A(EX_DW01_add_1__n125), .B(EX_DW01_add_1__n21), .C(EX_DW01_add_1__n333), .Y(EX_DW01_add_1__n652) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U411 ( .A(EX_DW01_add_1__n642), .Y(EX_DW01_add_1__n171) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U412 ( .A(EX_DW01_add_1__n597), .Y(EX_DW01_add_1__n172) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U413 ( .A(EX_DW01_add_1__n264), .Y(EX_DW01_add_1__n589) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U414 ( .A(EX_DW01_add_1__n584), .Y(EX_DW01_add_1__n173) );
  AO21x1_ASAP7_75t_R EX_DW01_add_1___U415 ( .A1(EX_DW01_add_1__n81), .A2(EX_DW01_add_1__n462), .B(EX_DW01_add_1__n350), .Y(EX_DW01_add_1__n508) );
  AO21x1_ASAP7_75t_R EX_DW01_add_1___U416 ( .A1(EX_DW01_add_1__n139), .A2(EX_DW01_add_1__n431), .B(EX_DW01_add_1__n497), .Y(EX_DW01_add_1__n493) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U417 ( .A(EX_DW01_add_1__n155), .Y(EX_DW01_add_1__n175) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U418 ( .A(EX_DW01_add_1__n629), .B(EX_DW01_add_1__n479), .Y(EX_DW01_add_1__n628) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U419 ( .A(EX_DW01_add_1__n177), .Y(EX_DW01_add_1__n176) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U420 ( .A(EX_DW01_add_1__n158), .Y(EX_DW01_add_1__n177) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U421 ( .A(EX_DW01_add_1__n163), .Y(EX_DW01_add_1__n178) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U422 ( .A(EX_DW01_add_1__n180), .Y(EX_DW01_add_1__n179) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U423 ( .A(EX_DW01_add_1__n166), .Y(EX_DW01_add_1__n180) );
  AO21x1_ASAP7_75t_R EX_DW01_add_1___U424 ( .A1(EX_DW01_add_1__n52), .A2(EX_DW01_add_1__n267), .B(EX_DW01_add_1__n428), .Y(EX_DW01_add_1__n596) );
  AO21x1_ASAP7_75t_R EX_DW01_add_1___U425 ( .A1(EX_DW01_add_1__n76), .A2(EX_DW01_add_1__n25), .B(EX_DW01_add_1__n237), .Y(EX_DW01_add_1__n570) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U426 ( .A(EX_DW01_add_1__n607), .Y(EX_DW01_add_1__n189) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U427 ( .A(EX_DW01_add_1__n183), .Y(EX_DW01_add_1__n182) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U428 ( .A(EX_DW01_add_1__n541), .Y(EX_DW01_add_1__n183) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U429 ( .A(EX_DW01_add_1__n498), .Y(EX_DW01_add_1__n184) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U430 ( .A(EX_DW01_add_1__n489), .Y(EX_DW01_add_1__n185) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U431 ( .A(EX_DW01_add_1__n571), .Y(EX_DW01_add_1__n186) );
  AO21x1_ASAP7_75t_R EX_DW01_add_1___U432 ( .A1(EX_DW01_add_1__n343), .A2(EX_DW01_add_1__n451), .B(EX_DW01_add_1__n637), .Y(EX_DW01_add_1__n635) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U433 ( .A(EX_DW01_add_1__n188), .Y(EX_DW01_add_1__n187) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U434 ( .A(EX_DW01_add_1__n157), .Y(EX_DW01_add_1__n188) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U435 ( .A(EX_DW01_add_1__n495), .B(EX_DW01_add_1__n427), .Y(EX_DW01_add_1__n494) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U436 ( .A(EX_DW01_add_1__n191), .Y(EX_DW01_add_1__n190) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U437 ( .A(EX_DW01_add_1__n528), .Y(EX_DW01_add_1__n191) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U438 ( .A(EX_DW01_add_1__n168), .Y(EX_DW01_add_1__n192) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U439 ( .A(EX_DW01_add_1__n236), .Y(EX_DW01_add_1__n193) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U440 ( .A(EX_DW01_add_1__n507), .Y(EX_DW01_add_1__n194) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U441 ( .A(EX_DW01_add_1__n587), .Y(EX_DW01_add_1__n195) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U442 ( .A(EX_DW01_add_1__n505), .Y(EX_DW01_add_1__n196) );
  AO21x1_ASAP7_75t_R EX_DW01_add_1___U443 ( .A1(EX_DW01_add_1__n21), .A2(EX_DW01_add_1__n22), .B(EX_DW01_add_1__n403), .Y(EX_DW01_add_1__n488) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U444 ( .A(EX_DW01_add_1__n198), .Y(EX_DW01_add_1__n197) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U445 ( .A(EX_DW01_add_1__n173), .Y(EX_DW01_add_1__n198) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U446 ( .A(EX_DW01_add_1__n585), .B(EX_DW01_add_1__n317), .Y(EX_DW01_add_1__n584) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U447 ( .A(EX_DW01_add_1__n200), .Y(EX_DW01_add_1__n199) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U448 ( .A(EX_DW01_add_1__n534), .Y(EX_DW01_add_1__n200) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U449 ( .A(EX_DW01_add_1__n202), .Y(EX_DW01_add_1__n201) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U450 ( .A(EX_DW01_add_1__n186), .Y(EX_DW01_add_1__n202) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U451 ( .A(EX_DW01_add_1__n204), .Y(EX_DW01_add_1__n203) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U452 ( .A(EX_DW01_add_1__n162), .Y(EX_DW01_add_1__n204) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U453 ( .A(EX_DW01_add_1__n486), .B(EX_DW01_add_1__n307), .Y(EX_DW01_add_1__n484) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U454 ( .A(EX_DW01_add_1__n161), .Y(EX_DW01_add_1__n206) );
  INVx6_ASAP7_75t_R EX_DW01_add_1___U455 ( .A(EX_DW01_add_1__n286), .Y(EX_DW01_add_1__n307) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U456 ( .A(EX_DW01_add_1__n455), .Y(EX_DW01_add_1__n614) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U457 ( .A(EX_DW01_add_1__n592), .Y(EX_DW01_add_1__n208) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U458 ( .A(EX_DW01_add_1__n604), .Y(EX_DW01_add_1__n209) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U459 ( .A(EX_DW01_add_1__n549), .Y(EX_DW01_add_1__n210) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U460 ( .A(EX_DW01_add_1__n212), .Y(EX_DW01_add_1__n211) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U461 ( .A(EX_DW01_add_1__n196), .Y(EX_DW01_add_1__n212) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U462 ( .A(EX_DW01_add_1__n477), .B(EX_DW01_add_1__n464), .Y(EX_DW01_add_1__n505) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U463 ( .A(EX_DW01_add_1__n214), .Y(EX_DW01_add_1__n213) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U464 ( .A(EX_DW01_add_1__n172), .Y(EX_DW01_add_1__n214) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U465 ( .A(EX_DW01_add_1__n589), .B(EX_DW01_add_1__n598), .Y(EX_DW01_add_1__n597) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U466 ( .A(EX_DW01_add_1__n216), .Y(EX_DW01_add_1__n215) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U467 ( .A(EX_DW01_add_1__n573), .Y(EX_DW01_add_1__n216) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U468 ( .A(EX_DW01_add_1__n197), .Y(EX_DW01_add_1__n217) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U469 ( .A(EX_DW01_add_1__n650), .Y(EX_DW01_add_1__n218) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U470 ( .A(EX_DW01_add_1__n564), .Y(EX_DW01_add_1__n219) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U471 ( .A(EX_DW01_add_1__n221), .Y(EX_DW01_add_1__n220) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U472 ( .A(EX_DW01_add_1__n208), .Y(EX_DW01_add_1__n221) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U473 ( .A(EX_DW01_add_1__n223), .Y(EX_DW01_add_1__n222) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U474 ( .A(EX_DW01_add_1__n170), .Y(EX_DW01_add_1__n223) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U475 ( .A(EX_DW01_add_1__n167), .Y(EX_DW01_add_1__n225) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U476 ( .A(EX_DW01_add_1__n169), .Y(EX_DW01_add_1__n227) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U477 ( .A(EX_DW01_add_1__n630), .Y(EX_DW01_add_1__n228) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U478 ( .A(EX_DW01_add_1__n195), .Y(EX_DW01_add_1__n230) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U479 ( .A(EX_DW01_add_1__n213), .Y(EX_DW01_add_1__n231) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U480 ( .A(EX_DW01_add_1__n187), .Y(EX_DW01_add_1__n232) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U481 ( .A(EX_DW01_add_1__n462), .B(EX_DW01_add_1__n448), .Y(EX_DW01_add_1__n522) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U482 ( .A(EX_DW01_add_1__n203), .Y(EX_DW01_add_1__n233) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U483 ( .A(EX_DW01_add_1__n184), .Y(EX_DW01_add_1__n234) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U484 ( .A(EX_DW01_add_1__n317), .B(EX_DW01_add_1__n375), .Y(EX_DW01_add_1__n236) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U485 ( .A(EX_DW01_add_1__n28), .B(EX_DW01_add_1__n450), .Y(EX_DW01_add_1__n573) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U486 ( .A(EX_DW01_add_1__n215), .Y(EX_DW01_add_1__n237) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U487 ( .A(EX_DW01_add_1__n657), .B(EX_DW01_add_1__n594), .Y(EX_DW01_add_1__n672) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U488 ( .A(EX_DW01_add_1__n159), .Y(EX_branch_addr[0]) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U489 ( .A(EX_DW01_add_1__n671), .Y(EX_branch_addr[1]) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U490 ( .A(EX_DW01_add_1__n626), .Y(EX_DW01_add_1__n251) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U491 ( .A(EX_DW01_add_1__n551), .Y(EX_DW01_add_1__n252) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U492 ( .A(EX_DW01_add_1__n662), .Y(EX_branch_addr[16]) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U493 ( .A(EX_DW01_add_1__n554), .Y(EX_DW01_add_1__n254) );
  AND4x1_ASAP7_75t_R EX_DW01_add_1___U494 ( .A(EX_DW01_add_1__n46), .B(EX_DW01_add_1__n48), .C(EX_DW01_add_1__n441), .D(EX_DW01_add_1__EX_DW01_add_1__n483), .Y(EX_DW01_add_1__n621) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U495 ( .A(EX_DW01_add_1__n563), .Y(EX_DW01_add_1__n255) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U496 ( .A(EX_DW01_add_1__n257), .Y(EX_DW01_add_1__n256) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U497 ( .A(EX_DW01_add_1__n575), .Y(EX_DW01_add_1__n257) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U498 ( .A(EX_DW01_add_1__n261), .Y(EX_DW01_add_1__n260) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U499 ( .A(EX_DW01_add_1__n254), .Y(EX_DW01_add_1__n261) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U500 ( .A(inst_addr[24]), .B(ID_EX_imm[24]), .Y(EX_DW01_add_1__n554) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U501 ( .A(EX_DW01_add_1__n566), .Y(EX_DW01_add_1__n263) );
  INVx3_ASAP7_75t_R EX_DW01_add_1___U502 ( .A(EX_DW01_add_1__n653), .Y(EX_DW01_add_1__n398) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U503 ( .A(EX_DW01_add_1__n562), .Y(EX_DW01_add_1__n415) );
  INVx6_ASAP7_75t_R EX_DW01_add_1___U504 ( .A(EX_DW01_add_1__n415), .Y(EX_DW01_add_1__n264) );
  AND4x1_ASAP7_75t_R EX_DW01_add_1___U505 ( .A(EX_DW01_add_1__n441), .B(EX_DW01_add_1__EX_DW01_add_1__n482), .C(EX_DW01_add_1__n48), .D(EX_DW01_add_1__EX_DW01_add_1__n483), .Y(EX_DW01_add_1__n561) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U506 ( .A(EX_DW01_add_1__n600), .Y(EX_DW01_add_1__n265) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U507 ( .A(EX_DW01_add_1__n419), .Y(EX_DW01_add_1__n266) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U508 ( .A(EX_DW01_add_1__n268), .Y(EX_DW01_add_1__n267) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U509 ( .A(EX_DW01_add_1__n270), .Y(EX_DW01_add_1__n269) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U510 ( .A(EX_DW01_add_1__n608), .Y(EX_DW01_add_1__n270) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U511 ( .A(EX_DW01_add_1__n276), .Y(EX_DW01_add_1__n275) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U512 ( .A(EX_DW01_add_1__n278), .Y(EX_DW01_add_1__n277) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U513 ( .A(EX_DW01_add_1__n543), .Y(EX_DW01_add_1__n278) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U514 ( .A(EX_DW01_add_1__n282), .Y(EX_DW01_add_1__n281) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U515 ( .A(EX_DW01_add_1__n256), .Y(EX_DW01_add_1__n282) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U516 ( .A(ID_EX_imm[22]), .B(inst_addr[22]), .Y(EX_DW01_add_1__n575) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U517 ( .A(inst_addr[12]), .B(ID_EX_imm[12]), .Y(EX_DW01_add_1__n626) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U518 ( .A(EX_DW01_add_1__n454), .Y(EX_DW01_add_1__n286) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U519 ( .A(EX_DW01_add_1__n288), .Y(EX_DW01_add_1__n287) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U520 ( .A(EX_DW01_add_1__n512), .Y(EX_DW01_add_1__n288) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U521 ( .A(EX_DW01_add_1__n290), .Y(EX_DW01_add_1__n289) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U522 ( .A(EX_DW01_add_1__n631), .Y(EX_DW01_add_1__n291) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U523 ( .A(EX_DW01_add_1__n633), .Y(EX_DW01_add_1__n292) );
  INVx6_ASAP7_75t_R EX_DW01_add_1___U524 ( .A(EX_DW01_add_1__n331), .Y(EX_DW01_add_1__n482) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U525 ( .A(EX_DW01_add_1__n457), .Y(EX_DW01_add_1__n295) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U526 ( .A(EX_DW01_add_1__n297), .Y(EX_DW01_add_1__n296) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U527 ( .A(EX_DW01_add_1__n538), .Y(EX_DW01_add_1__n297) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U528 ( .A(EX_DW01_add_1__n514), .Y(EX_DW01_add_1__n301) );
  AND2x6_ASAP7_75t_R EX_DW01_add_1___U529 ( .A(ID_EX_imm[19]), .B(inst_addr[19]), .Y(EX_DW01_add_1__n562) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U530 ( .A(EX_DW01_add_1__n520), .Y(EX_DW01_add_1__n303) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U531 ( .A(EX_DW01_add_1__n479), .B(EX_DW01_add_1__n70), .Y(EX_DW01_add_1__n560) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U532 ( .A(EX_DW01_add_1__n308), .Y(EX_DW01_add_1__n454) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U533 ( .A(EX_DW01_add_1__n310), .Y(EX_DW01_add_1__n309) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U534 ( .A(EX_DW01_add_1__n523), .Y(EX_DW01_add_1__n310) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U535 ( .A(EX_DW01_add_1__n526), .Y(EX_DW01_add_1__n524) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U536 ( .A(EX_DW01_add_1__n312), .Y(EX_DW01_add_1__n311) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U537 ( .A(EX_DW01_add_1__n531), .Y(EX_DW01_add_1__n312) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U538 ( .A(inst_addr[31]), .Y(EX_DW01_add_1__n314) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U539 ( .A(EX_DW01_add_1__n318), .Y(EX_DW01_add_1__n316) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U540 ( .A(EX_DW01_add_1__n318), .Y(EX_DW01_add_1__n317) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U541 ( .A(EX_DW01_add_1__n266), .Y(EX_DW01_add_1__n318) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U542 ( .A(ID_EX_imm[21]), .B(n2), .Y(EX_DW01_add_1__n419) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U543 ( .A(EX_DW01_add_1__n567), .Y(EX_DW01_add_1__n321) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U544 ( .A(inst_addr[1]), .B(ID_EX_imm[1]), .Y(EX_DW01_add_1__n653) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U545 ( .A(EX_DW01_add_1__n324), .Y(EX_DW01_add_1__n323) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U546 ( .A(EX_DW01_add_1__n506), .Y(EX_DW01_add_1__n324) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U547 ( .A(EX_DW01_add_1__n323), .Y(EX_DW01_add_1__n371) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U548 ( .A(ID_EX_imm[4]), .B(inst_addr[4]), .Y(EX_DW01_add_1__n506) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U549 ( .A(ID_EX_imm[25]), .B(n1), .Y(EX_DW01_add_1__n543) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U550 ( .A(EX_DW01_add_1__n328), .Y(EX_DW01_add_1__n327) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U551 ( .A(EX_DW01_add_1__n296), .Y(EX_DW01_add_1__n328) );
  INVx3_ASAP7_75t_R EX_DW01_add_1___U552 ( .A(EX_DW01_add_1__n327), .Y(EX_DW01_add_1__n449) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U553 ( .A(n4), .B(n786), .Y(EX_DW01_add_1__n602) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U554 ( .A(EX_DW01_add_1__n340), .Y(EX_DW01_add_1__n580) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U555 ( .A(EX_DW01_add_1__n260), .Y(EX_DW01_add_1__n330) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U556 ( .A(EX_DW01_add_1__n622), .Y(EX_DW01_add_1__n331) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U557 ( .A(EX_DW01_add_1__n510), .Y(EX_DW01_add_1__n437) );
  INVx6_ASAP7_75t_R EX_DW01_add_1___U558 ( .A(EX_DW01_add_1__n437), .Y(EX_DW01_add_1__n332) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U559 ( .A(EX_DW01_add_1__n591), .Y(EX_DW01_add_1__n334) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U560 ( .A(EX_DW01_add_1__n334), .Y(EX_DW01_add_1__n598) );
  OR2x6_ASAP7_75t_R EX_DW01_add_1___U561 ( .A(inst_addr[19]), .B(ID_EX_imm[19]), .Y(EX_DW01_add_1__n591) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U562 ( .A(EX_DW01_add_1__n569), .Y(EX_DW01_add_1__n335) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U563 ( .A(EX_DW01_add_1__n338), .Y(EX_DW01_add_1__n337) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U564 ( .A(EX_DW01_add_1__n649), .Y(EX_DW01_add_1__n338) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U565 ( .A(EX_DW01_add_1__n379), .B(EX_DW01_add_1__n339), .Y(EX_DW01_add_1__n650) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U566 ( .A(EX_DW01_add_1__n340), .Y(EX_DW01_add_1__n585) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U567 ( .A(EX_DW01_add_1__n342), .Y(EX_DW01_add_1__n341) );
  OA21x2_ASAP7_75t_R EX_DW01_add_1___U568 ( .A1(EX_DW01_add_1__n638), .A2(EX_DW01_add_1__n616), .B(EX_DW01_add_1__n283), .Y(EX_DW01_add_1__n343) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U569 ( .A(EX_DW01_add_1__n547), .Y(EX_DW01_add_1__n345) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U570 ( .A(EX_DW01_add_1__n335), .Y(EX_DW01_add_1__n347) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U571 ( .A(inst_addr[23]), .B(ID_EX_imm[23]), .Y(EX_DW01_add_1__n569) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U572 ( .A(inst_addr[17]), .B(ID_EX_imm[17]), .Y(EX_DW01_add_1__n610) );
  INVx3_ASAP7_75t_R EX_DW01_add_1___U573 ( .A(EX_DW01_add_1__n40), .Y(EX_DW01_add_1__n477) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U574 ( .A(EX_DW01_add_1__n309), .Y(EX_DW01_add_1__n350) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U575 ( .A(EX_DW01_add_1__n309), .Y(EX_DW01_add_1__n448) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U576 ( .A(EX_DW01_add_1__n582), .B(EX_DW01_add_1__n466), .Y(EX_DW01_add_1__n587) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U577 ( .A(EX_DW01_add_1__n511), .Y(EX_DW01_add_1__n396) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U578 ( .A(EX_DW01_add_1__n535), .B(EX_DW01_add_1__n92), .Y(EX_DW01_add_1__n541) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U579 ( .A(EX_DW01_add_1__n182), .Y(EX_DW01_add_1__n355) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U580 ( .A(EX_DW01_add_1__n658), .Y(EX_DW01_add_1__n356) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U581 ( .A(EX_DW01_add_1__n360), .Y(EX_DW01_add_1__n359) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U582 ( .A(EX_DW01_add_1__n171), .Y(EX_DW01_add_1__n360) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U583 ( .A(EX_DW01_add_1__n482), .Y(EX_DW01_add_1__n637) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U584 ( .A(EX_DW01_add_1__n209), .Y(EX_DW01_add_1__n362) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U585 ( .A(EX_DW01_add_1__n364), .Y(EX_DW01_add_1__n363) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U586 ( .A(EX_DW01_add_1__n185), .Y(EX_DW01_add_1__n364) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U587 ( .A(EX_DW01_add_1__n333), .Y(EX_DW01_add_1__n490) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U588 ( .A(EX_DW01_add_1__n593), .B(EX_DW01_add_1__n398), .Y(EX_DW01_add_1__n592) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U589 ( .A(EX_DW01_add_1__n220), .Y(EX_DW01_add_1__n365) );
  XOR2x2_ASAP7_75t_R EX_DW01_add_1___U590 ( .A(EX_DW01_add_1__n526), .B(EX_DW01_add_1__n365), .Y(EX_DW01_add_1__n671) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U591 ( .A(EX_DW01_add_1__n613), .B(EX_DW01_add_1__n472), .Y(EX_DW01_add_1__n612) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U592 ( .A(EX_DW01_add_1__n578), .B(EX_DW01_add_1__n579), .Y(EX_DW01_add_1__n577) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U593 ( .A(EX_DW01_add_1__n176), .Y(EX_DW01_add_1__n367) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U594 ( .A(EX_DW01_add_1__n321), .Y(EX_DW01_add_1__n368) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U595 ( .A(EX_DW01_add_1__n609), .B(EX_DW01_add_1__n455), .Y(EX_DW01_add_1__n615) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U596 ( .A(EX_DW01_add_1__n179), .Y(EX_DW01_add_1__n369) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U597 ( .A(EX_DW01_add_1__n429), .B(EX_DW01_add_1__n625), .Y(EX_DW01_add_1__n648) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U598 ( .A(EX_DW01_add_1__n371), .Y(EX_DW01_add_1__n504) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U599 ( .A(EX_DW01_add_1__n301), .Y(EX_DW01_add_1__n373) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U600 ( .A(EX_DW01_add_1__n580), .B(EX_DW01_add_1__n376), .Y(EX_DW01_add_1__n574) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U601 ( .A(EX_DW01_add_1__n410), .Y(EX_DW01_add_1__n376) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U602 ( .A(EX_DW01_add_1__n402), .B(EX_DW01_add_1__n378), .Y(EX_DW01_add_1__n631) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U603 ( .A(EX_DW01_add_1__n291), .Y(EX_DW01_add_1__n377) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U604 ( .A(EX_DW01_add_1__n465), .B(EX_DW01_add_1__n482), .Y(EX_DW01_add_1__n633) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U605 ( .A(EX_DW01_add_1__n292), .Y(EX_DW01_add_1__n378) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U606 ( .A(EX_DW01_add_1__n255), .Y(EX_DW01_add_1__n380) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U607 ( .A(EX_DW01_add_1__n497), .B(EX_DW01_add_1__n427), .Y(EX_DW01_add_1__n656) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U608 ( .A(EX_DW01_add_1__n502), .B(EX_DW01_add_1__n477), .Y(EX_DW01_add_1__n654) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U609 ( .A(EX_DW01_add_1__n454), .B(EX_DW01_add_1__n289), .Y(EX_DW01_add_1__n644) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U610 ( .A(EX_DW01_add_1__n645), .Y(EX_DW01_add_1__n384) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U611 ( .A(EX_DW01_add_1__n386), .Y(EX_DW01_add_1__n385) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U612 ( .A(EX_DW01_add_1__n356), .Y(EX_DW01_add_1__n386) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U613 ( .A(EX_DW01_add_1__n385), .Y(EX_DW01_add_1__n594) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U614 ( .A(EX_DW01_add_1__n388), .Y(EX_DW01_add_1__n387) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U615 ( .A(EX_DW01_add_1__n219), .Y(EX_DW01_add_1__n388) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U616 ( .A(EX_DW01_add_1__n545), .Y(EX_DW01_add_1__n389) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U617 ( .A(EX_DW01_add_1__n391), .Y(EX_DW01_add_1__n390) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U618 ( .A(EX_DW01_add_1__n303), .Y(EX_DW01_add_1__n391) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U619 ( .A(EX_DW01_add_1__n289), .B(EX_DW01_add_1__n490), .Y(EX_DW01_add_1__n489) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U620 ( .A(EX_DW01_add_1__n363), .Y(EX_DW01_add_1__n392) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U621 ( .A(EX_DW01_add_1__n486), .Y(EX_DW01_add_1__n651) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U622 ( .A(EX_DW01_add_1__n651), .Y(EX_DW01_add_1__n397) );
  AND2x4_ASAP7_75t_R EX_DW01_add_1___U623 ( .A(n786), .B(n4), .Y(EX_DW01_add_1__n600) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U624 ( .A(EX_DW01_add_1__n401), .Y(EX_DW01_add_1__n400) );
  BUFx12f_ASAP7_75t_R EX_DW01_add_1___U625 ( .A(EX_DW01_add_1__n496), .Y(EX_DW01_add_1__n401) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U626 ( .A(EX_DW01_add_1__n425), .Y(EX_DW01_add_1__n403) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U627 ( .A(EX_DW01_add_1__n518), .Y(EX_DW01_add_1__n405) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U628 ( .A(EX_DW01_add_1__n637), .B(EX_DW01_add_1__n643), .Y(EX_DW01_add_1__n642) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U629 ( .A(EX_DW01_add_1__n359), .Y(EX_DW01_add_1__n406) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U630 ( .A(EX_DW01_add_1__n380), .B(EX_DW01_add_1__n329), .Y(EX_DW01_add_1__n564) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U631 ( .A(EX_DW01_add_1__n387), .Y(EX_DW01_add_1__n409) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U632 ( .A(EX_DW01_add_1__n305), .Y(EX_DW01_add_1__n466) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U633 ( .A(EX_DW01_add_1__n421), .Y(EX_DW01_add_1__n420) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U634 ( .A(EX_DW01_add_1__n210), .Y(EX_DW01_add_1__n421) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U635 ( .A(EX_DW01_add_1__n164), .Y(EX_DW01_add_1__n424) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U636 ( .A(EX_DW01_add_1__n521), .B(EX_DW01_add_1__n390), .Y(EX_DW01_add_1__n515) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U637 ( .A(EX_DW01_add_1__n384), .Y(EX_DW01_add_1__n429) );
  INVx6_ASAP7_75t_R EX_DW01_add_1___U638 ( .A(EX_DW01_add_1__n389), .Y(EX_DW01_add_1__n430) );
  INVx3_ASAP7_75t_R EX_DW01_add_1___U639 ( .A(EX_DW01_add_1__n430), .Y(EX_DW01_add_1__n535) );
  OA21x2_ASAP7_75t_R EX_DW01_add_1___U640 ( .A1(EX_DW01_add_1__n434), .A2(EX_DW01_add_1__n130), .B(EX_DW01_add_1__n433), .Y(EX_DW01_add_1__n519) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U641 ( .A(ID_EX_imm[28]), .B(inst_addr[28]), .Y(EX_DW01_add_1__n531) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U642 ( .A(EX_DW01_add_1__n311), .Y(EX_DW01_add_1__n433) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U643 ( .A(EX_DW01_add_1__n529), .Y(EX_DW01_add_1__n434) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U644 ( .A(EX_DW01_add_1__n211), .Y(EX_DW01_add_1__n442) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U645 ( .A(EX_DW01_add_1__n572), .B(EX_DW01_add_1__n11), .Y(EX_DW01_add_1__n571) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U646 ( .A(EX_DW01_add_1__n201), .Y(EX_DW01_add_1__n443) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U647 ( .A(EX_DW01_add_1__n402), .B(EX_DW01_add_1__n465), .Y(EX_DW01_add_1__n636) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U648 ( .A(EX_DW01_add_1__n222), .Y(EX_DW01_add_1__n444) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U649 ( .A(inst_addr[10]), .B(ID_EX_imm[10]), .Y(EX_DW01_add_1__n649) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U650 ( .A(ID_EX_imm[27]), .B(inst_addr[27]), .Y(EX_DW01_add_1__n538) );
  XNOR2x2_ASAP7_75t_R EX_DW01_add_1___U651 ( .A(ID_EX_imm[31]), .B(EX_DW01_add_1__n314), .Y(EX_DW01_add_1__n512) );
  INVx4_ASAP7_75t_R EX_DW01_add_1___U652 ( .A(EX_DW01_add_1__n263), .Y(EX_DW01_add_1__n450) );
  AND2x2_ASAP7_75t_R EX_DW01_add_1___U653 ( .A(ID_EX_imm[16]), .B(inst_addr[16]), .Y(EX_DW01_add_1__n607) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U654 ( .A(EX_DW01_add_1__n606), .Y(EX_DW01_add_1__n456) );
  BUFx4f_ASAP7_75t_R EX_DW01_add_1___U655 ( .A(EX_DW01_add_1__n458), .Y(EX_DW01_add_1__n457) );
  BUFx3_ASAP7_75t_R EX_DW01_add_1___U656 ( .A(EX_DW01_add_1__n294), .Y(EX_DW01_add_1__n458) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U657 ( .A(EX_DW01_add_1__n460), .B(EX_DW01_add_1__n548), .Y(EX_DW01_add_1__n549) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U658 ( .A(EX_DW01_add_1__n420), .Y(EX_DW01_add_1__n459) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U659 ( .A(EX_DW01_add_1__n326), .Y(EX_DW01_add_1__n550) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U660 ( .A(EX_DW01_add_1__n550), .Y(EX_DW01_add_1__n460) );
  INVx2_ASAP7_75t_R EX_DW01_add_1___U661 ( .A(EX_DW01_add_1__n407), .Y(EX_DW01_add_1__n548) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U662 ( .A(EX_DW01_add_1__n463), .Y(EX_DW01_add_1__n462) );
  BUFx6f_ASAP7_75t_R EX_DW01_add_1___U663 ( .A(EX_DW01_add_1__n353), .Y(EX_DW01_add_1__n634) );
  INVx3_ASAP7_75t_R EX_DW01_add_1___U664 ( .A(EX_DW01_add_1__n634), .Y(EX_DW01_add_1__n465) );
  OA21x2_ASAP7_75t_R EX_DW01_add_1___U665 ( .A1(EX_DW01_add_1__n13), .A2(EX_DW01_add_1__n264), .B(EX_DW01_add_1__n380), .Y(EX_DW01_add_1__n551) );
  OA21x2_ASAP7_75t_R EX_DW01_add_1___U666 ( .A1(EX_DW01_add_1__n93), .A2(EX_DW01_add_1__n150), .B(EX_DW01_add_1__n126), .Y(EX_DW01_add_1__n552) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U667 ( .A(EX_DW01_add_1__n470), .B(EX_DW01_add_1__n352), .Y(EX_DW01_add_1__n604) );
  BUFx2_ASAP7_75t_R EX_DW01_add_1___U668 ( .A(EX_DW01_add_1__n399), .Y(EX_DW01_add_1__n605) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U669 ( .A(EX_DW01_add_1__n605), .Y(EX_DW01_add_1__n470) );
  INVx3_ASAP7_75t_R EX_DW01_add_1___U670 ( .A(EX_DW01_add_1__n500), .Y(EX_DW01_add_1__n473) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U671 ( .A(EX_DW01_add_1__n589), .B(EX_DW01_add_1__n315), .Y(EX_DW01_add_1__n588) );
  XOR2x2_ASAP7_75t_R EX_DW01_add_1___U672 ( .A(ID_EX_imm[29]), .B(inst_addr[29]), .Y(EX_DW01_add_1__n528) );
  XOR2x2_ASAP7_75t_R EX_DW01_add_1___U673 ( .A(ID_EX_imm[30]), .B(inst_addr[30]), .Y(EX_DW01_add_1__n518) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U674 ( .A(inst_addr[30]), .B(ID_EX_imm[30]), .Y(EX_DW01_add_1__n514) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U675 ( .A(inst_addr[29]), .B(ID_EX_imm[29]), .Y(EX_DW01_add_1__n520) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U676 ( .A(inst_addr[28]), .B(ID_EX_imm[28]), .Y(EX_DW01_add_1__n532) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U677 ( .A(inst_addr[27]), .B(ID_EX_imm[27]), .Y(EX_DW01_add_1__n536) );
  AOI311xp33_ASAP7_75t_R EX_DW01_add_1___U678 ( .A1(EX_DW01_add_1__n100), .A2(EX_DW01_add_1__n135), .A3(EX_DW01_add_1__n332), .B(EX_DW01_add_1__n54), .C(
        n481), .Y(EX_DW01_add_1__n556) );
  A2O1A1Ixp33_ASAP7_75t_R EX_DW01_add_1___U679 ( .A1(EX_DW01_add_1__n28), .A2(EX_DW01_add_1__n450), .B(EX_DW01_add_1__n11), .C(EX_DW01_add_1__n368), .Y(
        n553) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U680 ( .A(EX_DW01_add_1__n368), .Y(EX_DW01_add_1__n572) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U681 ( .A(EX_DW01_add_1__n450), .Y(EX_DW01_add_1__n579) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U682 ( .A(EX_DW01_add_1__n281), .Y(EX_DW01_add_1__n578) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U683 ( .A(inst_addr[20]), .B(ID_EX_imm[20]), .Y(EX_DW01_add_1__n582) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U684 ( .A(EX_DW01_add_1__n298), .Y(EX_DW01_add_1__n593) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U685 ( .A(EX_DW01_add_1__n414), .Y(EX_DW01_add_1__n613) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U686 ( .A(ID_EX_imm[16]), .B(EX_DW01_add_1__n69), .Y(EX_DW01_add_1__n609) );
  INVx1_ASAP7_75t_R EX_DW01_add_1___U687 ( .A(EX_DW01_add_1__n283), .Y(EX_DW01_add_1__n643) );
  A2O1A1Ixp33_ASAP7_75t_R EX_DW01_add_1___U688 ( .A1(EX_DW01_add_1__n259), .A2(EX_DW01_add_1__n468), .B(EX_DW01_add_1__n481), .C(EX_DW01_add_1__n436), .Y(
        n641) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U689 ( .A(inst_addr[2]), .B(ID_EX_imm[2]), .Y(EX_DW01_add_1__n509) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U690 ( .A(inst_addr[3]), .B(n762), .Y(EX_DW01_add_1__n511) );
  OR2x2_ASAP7_75t_R EX_DW01_add_1___U691 ( .A(inst_addr[0]), .B(n731), .Y(EX_DW01_add_1__n658) );



  BUFx5_ASAP7_75t_R EX___U1 ( .A(ID_EX_inst_addr[25]), .Y(EX__n1) );
  BUFx12f_ASAP7_75t_R EX___U2 ( .A(ID_EX_inst_addr[21]), .Y(EX__n2) );
  BUFx12f_ASAP7_75t_R EX___U3 ( .A(ID_EX_inst_addr[18]), .Y(EX__n4) );
  BUFx24_ASAP7_75t_R EX___U4 ( .A(EX__n1290), .Y(EX__n1281) );
  BUFx24_ASAP7_75t_R EX___U5 ( .A(EX__n1290), .Y(EX__n1282) );
  BUFx24_ASAP7_75t_R EX___U6 ( .A(EX__n1290), .Y(EX__n1283) );
  INVx1_ASAP7_75t_R EX___U7 ( .A(EX__n1202), .Y(EX_read_reg_data_2[11]) );
  BUFx2_ASAP7_75t_R EX___U8 ( .A(EX__n533), .Y(EX__n532) );
  HB1xp67_ASAP7_75t_R EX___U9 ( .A(EX__ALU_zero), .Y(EX__n5) );
  BUFx2_ASAP7_75t_R EX___U10 ( .A(EX__n512), .Y(EX__n831) );
  HB1xp67_ASAP7_75t_R EX___U11 ( .A(EX__n1617), .Y(EX__n512) );
  AOI21xp5_ASAP7_75t_R EX___U12 ( .A1(EX__n32), .A2(EX__n1569), .B(EX__EX__n692), .Y(EX__n6) );
  AOI21xp5_ASAP7_75t_R EX___U13 ( .A1(EX__n7), .A2(forwarding_MEM_WB[13]), .B(EX__n646), 
        .Y(EX__n1630) );
  CKINVDCx20_ASAP7_75t_R EX___U14 ( .A(EX__n1283), .Y(EX__n7) );
  INVxp67_ASAP7_75t_R EX___U15 ( .A(forwarding_MEM_WB[13]), .Y(EX__n41) );
  HB1xp67_ASAP7_75t_R EX___U16 ( .A(EX__n905), .Y(EX__n904) );
  INVxp67_ASAP7_75t_R EX___U17 ( .A(EX__n904), .Y(EX_read_reg_data_2[21]) );
  HB1xp67_ASAP7_75t_R EX___U18 ( .A(n56), .Y(EX__n8) );
  HB1xp67_ASAP7_75t_R EX___U19 ( .A(EX__n405), .Y(EX__n533) );
  BUFx2_ASAP7_75t_R EX___U20 ( .A(EX__n721), .Y(EX__n1202) );
  HB1xp67_ASAP7_75t_R EX___U21 ( .A(EX__n722), .Y(EX__n721) );
  HB1xp67_ASAP7_75t_R EX___U22 ( .A(ID_EX_imm[13]), .Y(EX__n1532) );
  HB1xp67_ASAP7_75t_R EX___U23 ( .A(EX__n531), .Y(EX__n722) );
  INVxp33_ASAP7_75t_R EX___U24 ( .A(ID_EX_imm[22]), .Y(EX__n1503) );
  HB1xp67_ASAP7_75t_R EX___U25 ( .A(EX_read_reg_data_2[2]), .Y(EX__n1567) );
  INVxp67_ASAP7_75t_R EX___U26 ( .A(EX__n1567), .Y(EX__n1254) );
  INVxp67_ASAP7_75t_R EX___U27 ( .A(EX__n576), .Y(EX_read_reg_data_2[2]) );
  HB1xp67_ASAP7_75t_R EX___U28 ( .A(EX__n577), .Y(EX__n576) );
  HB1xp67_ASAP7_75t_R EX___U29 ( .A(EX__n1635), .Y(EX__n405) );
  AOI21xp5_ASAP7_75t_R EX___U30 ( .A1(EX__n37), .A2(forwarding_MEM_WB[8]), .B(EX__n534), 
        .Y(EX__n1635) );
  HB1xp67_ASAP7_75t_R EX___U31 ( .A(forwarding_MEM_WB[1]), .Y(EX__n1569) );
  HB1xp67_ASAP7_75t_R EX___U32 ( .A(EX__n1632), .Y(EX__n531) );
  HB1xp67_ASAP7_75t_R EX___U33 ( .A(EX__n18), .Y(EX__n577) );
  INVxp67_ASAP7_75t_R EX___U34 ( .A(EX__n1621), .Y(EX_read_reg_data_2[22]) );
  AOI21xp5_ASAP7_75t_R EX___U35 ( .A1(forwarding_MEM_WB[22]), .A2(EX__n43), .B(EX__n681), 
        .Y(EX__n1621) );
  INVxp67_ASAP7_75t_R EX___U36 ( .A(EX__n834), .Y(EX_read_reg_data_2[20]) );
  BUFx2_ASAP7_75t_R EX___U37 ( .A(EX_read_reg_data_2[28]), .Y(EX__n1483) );
  HB1xp67_ASAP7_75t_R EX___U38 ( .A(EX__n835), .Y(EX__n834) );
  HB1xp67_ASAP7_75t_R EX___U39 ( .A(ID_EX_inst_addr[1]), .Y(EX__n10) );
  HB1xp67_ASAP7_75t_R EX___U40 ( .A(ID_EX_imm[9]), .Y(EX__n1544) );
  BUFx2_ASAP7_75t_R EX___U41 ( .A(EX__n825), .Y(EX__n823) );
  HB1xp67_ASAP7_75t_R EX___U42 ( .A(EX__n1481), .Y(EX__n825) );
  AOI21x1_ASAP7_75t_R EX___U43 ( .A1(EX__n11), .A2(forwarding_MEM_WB[27]), .B(EX__n718), 
        .Y(EX__n1616) );
  CKINVDCx20_ASAP7_75t_R EX___U44 ( .A(EX__n1287), .Y(EX__n11) );
  HB1xp67_ASAP7_75t_R EX___U45 ( .A(EX__n1623), .Y(EX__n835) );
  INVxp33_ASAP7_75t_R EX___U46 ( .A(EX__n46), .Y(EX__n1623) );
  INVxp33_ASAP7_75t_R EX___U47 ( .A(ID_EX_imm[6]), .Y(EX__n1556) );
  BUFx3_ASAP7_75t_R EX___U48 ( .A(ID_EX_imm[0]), .Y(EX__n731) );
  HB1xp67_ASAP7_75t_R EX___U49 ( .A(ID_EX_inst_addr[27]), .Y(EX__n12) );
  INVx1_ASAP7_75t_R EX___U50 ( .A(forwarding_MEM_WB[30]), .Y(EX__n13) );
  INVxp33_ASAP7_75t_R EX___U51 ( .A(EX__n13), .Y(EX__n14) );
  HB1xp67_ASAP7_75t_R EX___U52 ( .A(ID_EX_inst_addr[9]), .Y(EX__n15) );
  HB1xp67_ASAP7_75t_R EX___U53 ( .A(ID_EX_inst_addr[12]), .Y(EX__n49) );
  AOI21xp5_ASAP7_75t_R EX___U54 ( .A1(EX__n16), .A2(forwarding_MEM_WB[11]), .B(EX__n723), 
        .Y(EX__EX__n1632) );
  CKINVDCx20_ASAP7_75t_R EX___U55 ( .A(EX__n1282), .Y(EX__n16) );
  HB1xp67_ASAP7_75t_R EX___U56 ( .A(ID_EX_inst_addr[13]), .Y(EX__n17) );
  AOI21xp5_ASAP7_75t_R EX___U57 ( .A1(forwarding_MEM_WB[2]), .A2(EX__n53), .B(EX__n54), .Y(
        n18) );
  INVxp67_ASAP7_75t_R EX___U58 ( .A(EX__n1084), .Y(EX__n805) );
  HB1xp67_ASAP7_75t_R EX___U59 ( .A(ID_EX_imm[12]), .Y(EX__n19) );
  HB1xp67_ASAP7_75t_R EX___U60 ( .A(ID_EX_inst_addr[28]), .Y(EX__n20) );
  BUFx2_ASAP7_75t_R EX___U61 ( .A(EX__n869), .Y(EX__n867) );
  HB1xp67_ASAP7_75t_R EX___U62 ( .A(forwarding_MEM_WB[3]), .Y(EX__n869) );
  HB1xp67_ASAP7_75t_R EX___U63 ( .A(ID_EX_inst_addr[10]), .Y(EX__n21) );
  HB1xp67_ASAP7_75t_R EX___U64 ( .A(ID_EX_inst_addr[5]), .Y(EX__n22) );
  INVx2_ASAP7_75t_R EX___U65 ( .A(EX__n914), .Y(EX__n557) );
  INVx2_ASAP7_75t_R EX___U66 ( .A(EX__n19), .Y(EX__n1535) );
  INVx2_ASAP7_75t_R EX___U67 ( .A(forwarding_MEM_WB[16]), .Y(EX__n733) );
  INVx2_ASAP7_75t_R EX___U68 ( .A(EX__n557), .Y(EX__n976) );
  HB1xp67_ASAP7_75t_R EX___U69 ( .A(n58), .Y(EX__n23) );
  HB1xp67_ASAP7_75t_R EX___U70 ( .A(ID_EX_inst_addr[6]), .Y(EX__n24) );
  INVxp33_ASAP7_75t_R EX___U71 ( .A(ID_EX_imm[28]), .Y(EX__n1482) );
  HB1xp67_ASAP7_75t_R EX___U72 ( .A(ID_EX_inst_addr[2]), .Y(EX__n25) );
  INVx1_ASAP7_75t_R EX___U73 ( .A(EX__n917), .Y(EX__n65) );
  INVx2_ASAP7_75t_R EX___U74 ( .A(forwarding_MEM_WB[24]), .Y(EX__n1133) );
  INVxp67_ASAP7_75t_R EX___U75 ( .A(EX__n1618), .Y(EX__n639) );
  BUFx2_ASAP7_75t_R EX___U76 ( .A(EX__n984), .Y(EX__n983) );
  INVxp67_ASAP7_75t_R EX___U77 ( .A(EX__n569), .Y(EX_read_reg_data_2[23]) );
  HB1xp67_ASAP7_75t_R EX___U78 ( .A(EX__n1620), .Y(EX__n569) );
  INVxp67_ASAP7_75t_R EX___U79 ( .A(forwarding_MEM_WB[15]), .Y(EX__n26) );
  HB1xp67_ASAP7_75t_R EX___U80 ( .A(EX__n1494), .Y(EX__n984) );
  INVxp67_ASAP7_75t_R EX___U81 ( .A(forwarding_MEM_WB[31]), .Y(EX__n785) );
  HB1xp67_ASAP7_75t_R EX___U82 ( .A(EX_read_reg_data_2[31]), .Y(EX__n1473) );
  INVx1_ASAP7_75t_R EX___U83 ( .A(EX__n1006), .Y(EX__n52) );
  HB1xp67_ASAP7_75t_R EX___U84 ( .A(EX__n639), .Y(EX__n1494) );
  INVx1_ASAP7_75t_R EX___U85 ( .A(EX__n855), .Y(EX__n54) );
  HB1xp67_ASAP7_75t_R EX___U86 ( .A(EX__n825), .Y(EX__n824) );
  INVxp67_ASAP7_75t_R EX___U87 ( .A(EX__n824), .Y(EX__n884) );
  BUFx2_ASAP7_75t_R EX___U88 ( .A(EX__n880), .Y(EX__n879) );
  HB1xp67_ASAP7_75t_R EX___U89 ( .A(EX__n985), .Y(EX__n897) );
  INVxp33_ASAP7_75t_R EX___U90 ( .A(EX__n1624), .Y(EX_read_reg_data_2[19]) );
  HB1xp67_ASAP7_75t_R EX___U91 ( .A(EX__n986), .Y(EX__n985) );
  INVxp67_ASAP7_75t_R EX___U92 ( .A(EX__n1497), .Y(EX__n1213) );
  HB1xp67_ASAP7_75t_R EX___U93 ( .A(ID_EX_imm[4]), .Y(EX__n434) );
  AOI21x1_ASAP7_75t_R EX___U94 ( .A1(EX__n44), .A2(forwarding_MEM_WB[25]), .B(EX__n1047), 
        .Y(EX__n1618) );
  BUFx2_ASAP7_75t_R EX___U95 ( .A(EX__n1039), .Y(EX__n1037) );
  HB1xp67_ASAP7_75t_R EX___U96 ( .A(forwarding_MEM_WB[19]), .Y(EX__n1039) );
  INVxp33_ASAP7_75t_R EX___U97 ( .A(ID_EX_imm[5]), .Y(EX__n1560) );
  HB1xp67_ASAP7_75t_R EX___U98 ( .A(ID_EX_inst_addr[4]), .Y(EX__n27) );
  HB1xp67_ASAP7_75t_R EX___U99 ( .A(forwarding_MEM_WB[23]), .Y(EX__n880) );
  HB1xp67_ASAP7_75t_R EX___U100 ( .A(EX__n671), .Y(EX__n986) );
  HB1xp67_ASAP7_75t_R EX___U101 ( .A(EX_read_reg_data_2[23]), .Y(EX__n1500) );
  INVxp67_ASAP7_75t_R EX___U102 ( .A(EX__n1500), .Y(EX__n1126) );
  HB1xp67_ASAP7_75t_R EX___U103 ( .A(forwarding_MEM_WB[10]), .Y(EX__n28) );
  INVx1_ASAP7_75t_R EX___U104 ( .A(forwarding_MEM_WB[10]), .Y(EX__n62) );
  HB1xp67_ASAP7_75t_R EX___U105 ( .A(EX__n731), .Y(EX__n29) );
  HB1xp67_ASAP7_75t_R EX___U106 ( .A(EX_read_reg_data_2[24]), .Y(EX__n1497) );
  INVx1_ASAP7_75t_R EX___U107 ( .A(forwarding_MEM_WB[21]), .Y(EX__n30) );
  HB1xp67_ASAP7_75t_R EX___U108 ( .A(ID_EX_imm[24]), .Y(EX__n1496) );
  BUFx3_ASAP7_75t_R EX___U109 ( .A(EX__n1000), .Y(EX_PCSrc) );
  INVxp33_ASAP7_75t_R EX___U110 ( .A(EX__n865), .Y(EX__n995) );
  HB1xp67_ASAP7_75t_R EX___U111 ( .A(EX_read_reg_data_2[21]), .Y(EX__n1508) );
  INVxp67_ASAP7_75t_R EX___U112 ( .A(EX__n1619), .Y(EX_read_reg_data_2[24]) );
  HB1xp67_ASAP7_75t_R EX___U113 ( .A(EX__n1624), .Y(EX__n671) );
  INVx1_ASAP7_75t_R EX___U114 ( .A(EX__n1637), .Y(EX_read_reg_data_2[5]) );
  INVx2_ASAP7_75t_R EX___U115 ( .A(EX__n1613), .Y(EX_read_reg_data_2[30]) );
  INVxp67_ASAP7_75t_R EX___U116 ( .A(EX__n1476), .Y(EX__n1168) );
  INVxp67_ASAP7_75t_R EX___U117 ( .A(EX__n939), .Y(EX__n1142) );
  HB1xp67_ASAP7_75t_R EX___U118 ( .A(EX__n940), .Y(EX__n939) );
  INVx2_ASAP7_75t_R EX___U119 ( .A(EX__n1628), .Y(EX_read_reg_data_2[15]) );
  INVxp67_ASAP7_75t_R EX___U120 ( .A(EX__n1527), .Y(EX__n1224) );
  HB1xp67_ASAP7_75t_R EX___U121 ( .A(EX__n404), .Y(EX__n905) );
  BUFx6f_ASAP7_75t_R EX___U122 ( .A(EX__n1506), .Y(EX__n865) );
  HB1xp67_ASAP7_75t_R EX___U123 ( .A(EX__n1622), .Y(EX__n404) );
  CKINVDCx20_ASAP7_75t_R EX___U124 ( .A(EX__n1288), .Y(EX__n32) );
  AO21x1_ASAP7_75t_R EX___U125 ( .A1(EX__n47), .A2(forwarding_MEM_WB[20]), .B(EX__n48), .Y(
        n46) );
  INVx1_ASAP7_75t_R EX___U126 ( .A(EX__n950), .Y(EX__n48) );
  HB1xp67_ASAP7_75t_R EX___U127 ( .A(EX__n14), .Y(EX__n866) );
  INVxp33_ASAP7_75t_R EX___U128 ( .A(EX__n1203), .Y(EX__n695) );
  BUFx3_ASAP7_75t_R EX___U129 ( .A(EX__n690), .Y(EX__n1203) );
  INVxp67_ASAP7_75t_R EX___U130 ( .A(forwarding_MEM_WB[12]), .Y(EX__n33) );
  INVxp33_ASAP7_75t_R EX___U131 ( .A(EX__n782), .Y(EX__n34) );
  INVxp67_ASAP7_75t_R EX___U132 ( .A(EX__n1146), .Y(EX_read_reg_data_2[12]) );
  HB1xp67_ASAP7_75t_R EX___U133 ( .A(EX__n935), .Y(EX__n1146) );
  INVxp67_ASAP7_75t_R EX___U134 ( .A(forwarding_MEM_WB[4]), .Y(EX__n35) );
  INVxp33_ASAP7_75t_R EX___U135 ( .A(EX__n822), .Y(EX__n36) );
  HB1xp67_ASAP7_75t_R EX___U136 ( .A(EX__n936), .Y(EX__n935) );
  CKINVDCx20_ASAP7_75t_R EX___U137 ( .A(EX__n1281), .Y(EX__n37) );
  HB1xp67_ASAP7_75t_R EX___U138 ( .A(EX__n35), .Y(EX__n822) );
  BUFx3_ASAP7_75t_R EX___U139 ( .A(ID_EX_inst_addr[3]), .Y(EX__n38) );
  HB1xp67_ASAP7_75t_R EX___U140 ( .A(ID_EX_imm[3]), .Y(EX__n763) );
  AO21x1_ASAP7_75t_R EX___U141 ( .A1(EX__n51), .A2(forwarding_MEM_WB[6]), .B(EX__n52), .Y(
        EX_read_reg_data_2[6]) );
  HB1xp67_ASAP7_75t_R EX___U142 ( .A(n39), .Y(EX__n39) );
  HB1xp67_ASAP7_75t_R EX___U143 ( .A(EX__n935), .Y(EX__n860) );
  HB1xp67_ASAP7_75t_R EX___U144 ( .A(EX__n34), .Y(EX__n1045) );
  BUFx2_ASAP7_75t_R EX___U145 ( .A(ID_EX_imm[3]), .Y(EX__n762) );
  HB1xp67_ASAP7_75t_R EX___U146 ( .A(ID_EX_imm[27]), .Y(EX__n40) );
  INVxp67_ASAP7_75t_R EX___U147 ( .A(forwarding_MEM_WB[7]), .Y(EX__n61) );
  HB1xp67_ASAP7_75t_R EX___U148 ( .A(EX__n1525), .Y(EX__n878) );
  BUFx6f_ASAP7_75t_R EX___U149 ( .A(EX__n1547), .Y(EX__n876) );
  INVxp67_ASAP7_75t_R EX___U150 ( .A(EX__n1614), .Y(EX_read_reg_data_2[29]) );
  HB1xp67_ASAP7_75t_R EX___U151 ( .A(forwarding_MEM_WB[31]), .Y(EX__n1471) );
  HB1xp67_ASAP7_75t_R EX___U152 ( .A(EX_read_reg_data_2[29]), .Y(EX__n1479) );
  INVxp67_ASAP7_75t_R EX___U153 ( .A(EX__n1479), .Y(EX__n1124) );
  BUFx3_ASAP7_75t_R EX___U154 ( .A(EX__n976), .Y(EX__n913) );
  HB1xp67_ASAP7_75t_R EX___U155 ( .A(EX_read_reg_data_2[15]), .Y(EX__n1527) );
  HB1xp67_ASAP7_75t_R EX___U156 ( .A(EX__n878), .Y(EX__n877) );
  BUFx3_ASAP7_75t_R EX___U157 ( .A(EX__n1627), .Y(EX__n914) );
  HB1xp67_ASAP7_75t_R EX___U158 ( .A(EX_read_reg_data_2[30]), .Y(EX__n1476) );
  BUFx2_ASAP7_75t_R EX___U159 ( .A(EX__n706), .Y(EX__n705) );
  HB1xp67_ASAP7_75t_R EX___U160 ( .A(EX__n410), .Y(EX__n706) );
  HB1xp67_ASAP7_75t_R EX___U161 ( .A(EX__n1612), .Y(EX__n410) );
  HB1xp67_ASAP7_75t_R EX___U162 ( .A(EX__n672), .Y(EX__n936) );
  INVx2_ASAP7_75t_R EX___U163 ( .A(EX__n656), .Y(EX_read_reg_data_2[7]) );
  BUFx3_ASAP7_75t_R EX___U164 ( .A(EX__n1636), .Y(EX__n656) );
  INVxp33_ASAP7_75t_R EX___U165 ( .A(EX__n41), .Y(EX__n42) );
  INVxp67_ASAP7_75t_R EX___U166 ( .A(EX__n521), .Y(EX__n943) );
  HB1xp67_ASAP7_75t_R EX___U167 ( .A(EX__n42), .Y(EX__n521) );
  CKINVDCx20_ASAP7_75t_R EX___U168 ( .A(EX__n1286), .Y(EX__n43) );
  CKINVDCx20_ASAP7_75t_R EX___U169 ( .A(EX__n624), .Y(EX__n44) );
  INVx1_ASAP7_75t_R EX___U170 ( .A(EX__n1154), .Y(EX_read_reg_data_2[25]) );
  HB1xp67_ASAP7_75t_R EX___U171 ( .A(EX__n1631), .Y(EX__n672) );
  HB1xp67_ASAP7_75t_R EX___U172 ( .A(EX__n33), .Y(EX__n782) );
  INVxp67_ASAP7_75t_R EX___U173 ( .A(EX__n1625), .Y(EX_read_reg_data_2[18]) );
  INVxp33_ASAP7_75t_R EX___U174 ( .A(EX__n709), .Y(EX__n911) );
  INVxp67_ASAP7_75t_R EX___U175 ( .A(EX__n1517), .Y(EX__n1221) );
  BUFx3_ASAP7_75t_R EX___U176 ( .A(EX__n1615), .Y(EX__n676) );
  CKINVDCx20_ASAP7_75t_R EX___U177 ( .A(EX__n1285), .Y(EX__n47) );
  BUFx3_ASAP7_75t_R EX___U178 ( .A(EX__n1639), .Y(EX__n673) );
  INVx2_ASAP7_75t_R EX___U179 ( .A(forwarding_MEM_WB[29]), .Y(EX__n989) );
  HB1xp67_ASAP7_75t_R EX___U180 ( .A(forwarding_MEM_WB[28]), .Y(EX__n1481) );
  CKINVDCx20_ASAP7_75t_R EX___U181 ( .A(EX__n1281), .Y(EX__n51) );
  CKINVDCx20_ASAP7_75t_R EX___U182 ( .A(EX__n1293), .Y(EX__n53) );
  HB1xp67_ASAP7_75t_R EX___U183 ( .A(EX__n869), .Y(EX__n868) );
  INVxp67_ASAP7_75t_R EX___U184 ( .A(EX__n1504), .Y(EX__n1163) );
  INVx1_ASAP7_75t_R EX___U185 ( .A(EX__n679), .Y(EX__n1050) );
  HB1xp67_ASAP7_75t_R EX___U186 ( .A(EX__n680), .Y(EX__n679) );
  BUFx3_ASAP7_75t_R EX___U187 ( .A(EX__n415), .Y(EX__n414) );
  HB1xp67_ASAP7_75t_R EX___U188 ( .A(EX__n982), .Y(EX__n981) );
  HB1xp67_ASAP7_75t_R EX___U189 ( .A(EX_read_reg_data_2[17]), .Y(EX__n1521) );
  INVx2_ASAP7_75t_R EX___U190 ( .A(EX__n823), .Y(EX__n883) );
  HB1xp67_ASAP7_75t_R EX___U191 ( .A(EX__n1565), .Y(EX__n944) );
  BUFx3_ASAP7_75t_R EX___U192 ( .A(EX__n573), .Y(EX__n572) );
  BUFx6f_ASAP7_75t_R EX___U193 ( .A(EX__n1519), .Y(EX__n982) );
  INVx2_ASAP7_75t_R EX___U194 ( .A(EX__n867), .Y(EX__n990) );
  AOI21x1_ASAP7_75t_R EX___U195 ( .A1(EX__n55), .A2(forwarding_MEM_WB[26]), .B(EX__n832), 
        .Y(EX__n1617) );
  CKINVDCx20_ASAP7_75t_R EX___U196 ( .A(EX__n1288), .Y(EX__n55) );
  BUFx3_ASAP7_75t_R EX___U197 ( .A(EX__n932), .Y(EX__n931) );
  BUFx3_ASAP7_75t_R EX___U198 ( .A(EX__n1626), .Y(EX__n826) );
  HB1xp67_ASAP7_75t_R EX___U199 ( .A(EX_read_reg_data_2[6]), .Y(EX__n729) );
  HB1xp67_ASAP7_75t_R EX___U200 ( .A(EX__n530), .Y(EX__n680) );
  HB1xp67_ASAP7_75t_R EX___U201 ( .A(EX__n1621), .Y(EX__n530) );
  INVxp33_ASAP7_75t_R EX___U202 ( .A(EX__n36), .Y(EX__n622) );
  AO22x1_ASAP7_75t_R EX___U203 ( .A1(EX__n434), .A2(ID_EX_ALUSrc), .B1(
        EX_read_reg_data_2[4]), .B2(EX__n1579), .Y(input_data_2[4]) );
  HB1xp67_ASAP7_75t_R EX___U204 ( .A(forwarding_MEM_WB[2]), .Y(EX__n1565) );
  HB1xp67_ASAP7_75t_R EX___U205 ( .A(EX__n1502), .Y(EX__n903) );
  HB1xp67_ASAP7_75t_R EX___U206 ( .A(ID_EX_imm[20]), .Y(EX__n56) );
  HB1xp67_ASAP7_75t_R EX___U207 ( .A(EX__n1555), .Y(EX__n842) );
  HB1xp67_ASAP7_75t_R EX___U208 ( .A(forwarding_MEM_WB[6]), .Y(EX__n1555) );
  INVxp33_ASAP7_75t_R EX___U209 ( .A(EX__n842), .Y(EX__n670) );
  INVx2_ASAP7_75t_R EX___U210 ( .A(forwarding_MEM_WB[17]), .Y(EX__n1043) );
  HB1xp67_ASAP7_75t_R EX___U211 ( .A(forwarding_MEM_WB[22]), .Y(EX__n1502) );
  INVx1_ASAP7_75t_R EX___U212 ( .A(EX__n1629), .Y(EX_read_reg_data_2[14]) );
  INVxp33_ASAP7_75t_R EX___U213 ( .A(EX__n838), .Y(EX__n1200) );
  HB1xp67_ASAP7_75t_R EX___U214 ( .A(EX__n874), .Y(EX__n873) );
  INVxp33_ASAP7_75t_R EX___U215 ( .A(EX__n944), .Y(EX__n804) );
  HB1xp67_ASAP7_75t_R EX___U216 ( .A(EX__n839), .Y(EX__n838) );
  HB1xp67_ASAP7_75t_R EX___U217 ( .A(EX__n1200), .Y(EX__n1530) );
  INVxp67_ASAP7_75t_R EX___U218 ( .A(EX__n1530), .Y(EX__n1172) );
  HB1xp67_ASAP7_75t_R EX___U219 ( .A(EX__n29), .Y(EX__n732) );
  HB1xp67_ASAP7_75t_R EX___U220 ( .A(ID_EX_inst_addr[22]), .Y(EX__n58) );
  HB1xp67_ASAP7_75t_R EX___U221 ( .A(EX__n40), .Y(EX__n1485) );
  INVx2_ASAP7_75t_R EX___U222 ( .A(forwarding_MEM_WB[9]), .Y(EX__n1040) );
  HB1xp67_ASAP7_75t_R EX___U223 ( .A(EX__n1569), .Y(EX__n945) );
  HB1xp67_ASAP7_75t_R EX___U224 ( .A(EX__n911), .Y(EX__n1517) );
  HB1xp67_ASAP7_75t_R EX___U225 ( .A(EX__n412), .Y(EX__n839) );
  HB1xp67_ASAP7_75t_R EX___U226 ( .A(EX__n1629), .Y(EX__n412) );
  BUFx6f_ASAP7_75t_R EX___U227 ( .A(forwarding_MEM_WB[14]), .Y(EX__n874) );
  HB1xp67_ASAP7_75t_R EX___U228 ( .A(EX__n710), .Y(EX__n709) );
  BUFx3_ASAP7_75t_R EX___U229 ( .A(EX__n1638), .Y(EX__n369) );
  INVxp33_ASAP7_75t_R EX___U230 ( .A(ID_EX_imm[8]), .Y(EX__n1548) );
  HB1xp67_ASAP7_75t_R EX___U231 ( .A(ID_EX_imm[15]), .Y(EX__n1526) );
  HB1xp67_ASAP7_75t_R EX___U232 ( .A(ID_EX_imm[10]), .Y(EX__n59) );
  INVxp33_ASAP7_75t_R EX___U234 ( .A(ID_EX_imm[26]), .Y(EX__n1489) );
  INVxp67_ASAP7_75t_R EX___U235 ( .A(EX__n902), .Y(EX__n1082) );
  HB1xp67_ASAP7_75t_R EX___U236 ( .A(EX__n1050), .Y(EX__n1504) );
  HB1xp67_ASAP7_75t_R EX___U237 ( .A(EX__n827), .Y(EX__n940) );
  HB1xp67_ASAP7_75t_R EX___U238 ( .A(EX__n1637), .Y(EX__n827) );
  INVx2_ASAP7_75t_R EX___U239 ( .A(EX__n872), .Y(EX__n997) );
  BUFx6f_ASAP7_75t_R EX___U240 ( .A(EX__n874), .Y(EX__n872) );
  HB1xp67_ASAP7_75t_R EX___U241 ( .A(EX__n903), .Y(EX__n902) );
  HB1xp67_ASAP7_75t_R EX___U242 ( .A(EX__n513), .Y(EX__n710) );
  HB1xp67_ASAP7_75t_R EX___U243 ( .A(EX__n1625), .Y(EX__n513) );
  INVx6_ASAP7_75t_R EX___U244 ( .A(EX__n584), .Y(EX__n882) );
  BUFx12f_ASAP7_75t_R EX___U245 ( .A(forwarding_MEM_WB[18]), .Y(EX__n584) );
  BUFx3_ASAP7_75t_R EX___U246 ( .A(EX__n1634), .Y(EX__n390) );
  AO21x1_ASAP7_75t_R EX___U247 ( .A1(EX__n64), .A2(forwarding_MEM_WB[0]), .B(EX__n65), .Y(
        n63) );
  INVxp67_ASAP7_75t_R EX___U248 ( .A(EX__n63), .Y(EX__n1640) );
  HB1xp67_ASAP7_75t_R EX___U249 ( .A(EX__n704), .Y(EX__n993) );
  INVxp33_ASAP7_75t_R EX___U250 ( .A(EX__n993), .Y(EX__n901) );
  INVxp33_ASAP7_75t_R EX___U251 ( .A(EX__n1202), .Y(EX__n726) );
  INVxp33_ASAP7_75t_R EX___U252 ( .A(forwarding_MEM_WB[27]), .Y(EX__n1042) );
  HB1xp67_ASAP7_75t_R EX___U253 ( .A(EX__n1559), .Y(EX__n704) );
  HB1xp67_ASAP7_75t_R EX___U254 ( .A(forwarding_MEM_WB[5]), .Y(EX__n1559) );
  HB1xp67_ASAP7_75t_R EX___U255 ( .A(forwarding_MEM_WB[11]), .Y(EX__n1084) );
  HB1xp67_ASAP7_75t_R EX___U256 ( .A(ID_EX_imm[1]), .Y(EX__n60) );
  HB1xp67_ASAP7_75t_R EX___U257 ( .A(EX__n60), .Y(EX__n1570) );
  HB1xp67_ASAP7_75t_R EX___U258 ( .A(forwarding_MEM_WB[15]), .Y(EX__n1525) );
  HB1xp67_ASAP7_75t_R EX___U259 ( .A(EX__n1039), .Y(EX__n1038) );
  INVxp67_ASAP7_75t_R EX___U260 ( .A(EX__n1561), .Y(EX__n1131) );
  HB1xp67_ASAP7_75t_R EX___U261 ( .A(EX__n1142), .Y(EX__n1561) );
  BUFx3_ASAP7_75t_R EX___U262 ( .A(EX__n717), .Y(EX__n716) );
  BUFx3_ASAP7_75t_R EX___U263 ( .A(EX__n1616), .Y(EX__n411) );
  INVxp33_ASAP7_75t_R EX___U264 ( .A(EX__n704), .Y(EX__n994) );
  HB1xp67_ASAP7_75t_R EX___U265 ( .A(EX__n901), .Y(EX__n863) );
  INVx2_ASAP7_75t_R EX___U266 ( .A(EX__n1037), .Y(EX__n1134) );
  HB1xp67_ASAP7_75t_R EX___U267 ( .A(EX__n1551), .Y(EX__n908) );
  HB1xp67_ASAP7_75t_R EX___U268 ( .A(forwarding_MEM_WB[7]), .Y(EX__n1551) );
  HB1xp67_ASAP7_75t_R EX___U269 ( .A(EX_read_reg_data_2[20]), .Y(EX__n1512) );
  HB1xp67_ASAP7_75t_R EX___U270 ( .A(EX_read_reg_data_2[10]), .Y(EX__n1542) );
  INVx2_ASAP7_75t_R EX___U271 ( .A(EX__n572), .Y(EX_read_reg_data_2[10]) );
  CKINVDCx20_ASAP7_75t_R EX___U272 ( .A(EX__n1085), .Y(EX__n64) );
  HB1xp67_ASAP7_75t_R EX___U273 ( .A(forwarding_MEM_WB[20]), .Y(EX__n1510) );
  HB1xp67_ASAP7_75t_R EX___U274 ( .A(EX__n1540), .Y(EX__n735) );
  HB1xp67_ASAP7_75t_R EX___U275 ( .A(EX__n871), .Y(EX__n870) );
  HB1xp67_ASAP7_75t_R EX___U276 ( .A(EX__n28), .Y(EX__n1540) );
  HB1xp67_ASAP7_75t_R EX___U277 ( .A(EX__n1510), .Y(EX__n1083) );
  HB1xp67_ASAP7_75t_R EX___U278 ( .A(EX_read_reg_data_2[0]), .Y(EX__n1577) );
  BUFx6f_ASAP7_75t_R EX___U279 ( .A(EX__n1574), .Y(EX__n871) );
  INVxp67_ASAP7_75t_R EX___U280 ( .A(EX__n580), .Y(EX_read_reg_data_2[0]) );
  HB1xp67_ASAP7_75t_R EX___U281 ( .A(EX__n581), .Y(EX__n580) );
  BUFx2_ASAP7_75t_R EX___U282 ( .A(ID_EX_imm[14]), .Y(EX__n1529) );
  BUFx3_ASAP7_75t_R EX___U283 ( .A(EX__n1633), .Y(EX__n413) );
  HB1xp67_ASAP7_75t_R EX___U284 ( .A(EX__n1640), .Y(EX__n581) );
  HB1xp67_ASAP7_75t_R EX___U285 ( .A(ID_EX_imm[2]), .Y(EX__n1566) );
  HB1xp67_ASAP7_75t_R EX___U286 ( .A(ID_EX_inst_addr[20]), .Y(EX__n67) );
  HB1xp67_ASAP7_75t_R EX___U287 ( .A(EX__n67), .Y(EX__n68) );
  INVxp33_ASAP7_75t_R EX___U288 ( .A(EX__n56), .Y(EX__n1511) );
  HB1xp67_ASAP7_75t_R EX___U289 ( .A(EX__n68), .Y(EX__n69) );
  HB1xp67_ASAP7_75t_R EX___U290 ( .A(EX__n59), .Y(EX__n730) );
  INVx2_ASAP7_75t_R EX___U291 ( .A(EX__n95), .Y(EX__n70) );
  BUFx2_ASAP7_75t_R EX___U292 ( .A(EX__n1299), .Y(EX__n71) );
  BUFx12f_ASAP7_75t_R EX___U293 ( .A(EX__n1299), .Y(EX__n72) );
  BUFx2_ASAP7_75t_R EX___U294 ( .A(EX__n1299), .Y(EX__n73) );
  BUFx2_ASAP7_75t_R EX___U295 ( .A(EX__n1299), .Y(EX__n74) );
  INVx2_ASAP7_75t_R EX___U296 ( .A(EX__n86), .Y(EX__n75) );
  CKINVDCx6p67_ASAP7_75t_R EX___U297 ( .A(ID_EX_ALUSrc), .Y(EX__n1579) );
  BUFx12f_ASAP7_75t_R EX___U298 ( .A(EX__n103), .Y(EX__n76) );
  BUFx12f_ASAP7_75t_R EX___U299 ( .A(EX__n103), .Y(EX__n77) );
  BUFx12f_ASAP7_75t_R EX___U300 ( .A(EX__n121), .Y(EX__n78) );
  BUFx12f_ASAP7_75t_R EX___U301 ( .A(EX__n121), .Y(EX__n79) );
  BUFx12f_ASAP7_75t_R EX___U302 ( .A(EX__n1304), .Y(EX__n80) );
  BUFx6f_ASAP7_75t_R EX___U303 ( .A(EX__n757), .Y(EX__n755) );
  INVx6_ASAP7_75t_R EX___U304 ( .A(EX__n105), .Y(EX__n104) );
  BUFx12f_ASAP7_75t_R EX___U305 ( .A(EX__n99), .Y(EX__n81) );
  BUFx3_ASAP7_75t_R EX___U306 ( .A(EX__n1356), .Y(EX__n82) );
  BUFx12f_ASAP7_75t_R EX___U307 ( .A(EX__n1356), .Y(EX__n83) );
  BUFx2_ASAP7_75t_R EX___U308 ( .A(EX__n1356), .Y(EX__n84) );
  BUFx2_ASAP7_75t_R EX___U309 ( .A(EX__n1356), .Y(EX__n85) );
  BUFx12f_ASAP7_75t_R EX___U310 ( .A(EX__n96), .Y(EX__n86) );
  BUFx12f_ASAP7_75t_R EX___U311 ( .A(EX__n96), .Y(EX__n87) );
  CKINVDCx20_ASAP7_75t_R EX___U312 ( .A(EX__n97), .Y(EX__n88) );
  BUFx12f_ASAP7_75t_R EX___U313 ( .A(EX__n926), .Y(EX__n105) );
  INVx6_ASAP7_75t_R EX___U314 ( .A(EX__n111), .Y(EX__n110) );
  BUFx2_ASAP7_75t_R EX___U315 ( .A(EX__n140), .Y(EX__n89) );
  BUFx12f_ASAP7_75t_R EX___U316 ( .A(EX__n91), .Y(EX__n90) );
  BUFx12f_ASAP7_75t_R EX___U317 ( .A(EX__n1343), .Y(EX__n91) );
  INVx6_ASAP7_75t_R EX___U318 ( .A(EX__n90), .Y(EX__n1205) );
  BUFx12f_ASAP7_75t_R EX___U319 ( .A(EX__n102), .Y(EX__n92) );
  BUFx12f_ASAP7_75t_R EX___U320 ( .A(EX__n102), .Y(EX__n93) );
  BUFx12f_ASAP7_75t_R EX___U321 ( .A(EX__n87), .Y(EX__n94) );
  BUFx12f_ASAP7_75t_R EX___U322 ( .A(EX__n86), .Y(EX__n95) );
  BUFx12f_ASAP7_75t_R EX___U323 ( .A(EX__n1317), .Y(EX__n96) );
  BUFx16f_ASAP7_75t_R EX___U324 ( .A(EX__n104), .Y(EX__n97) );
  CKINVDCx20_ASAP7_75t_R EX___U325 ( .A(EX__n106), .Y(EX__n98) );
  BUFx12f_ASAP7_75t_R EX___U326 ( .A(EX__n970), .Y(EX__n111) );
  BUFx12f_ASAP7_75t_R EX___U327 ( .A(EX__n885), .Y(EX__n99) );
  CKINVDCx9p33_ASAP7_75t_R EX___U328 ( .A(EX__n113), .Y(EX__n148) );
  BUFx12f_ASAP7_75t_R EX___U329 ( .A(EX__n93), .Y(EX__n100) );
  BUFx12f_ASAP7_75t_R EX___U330 ( .A(EX__n92), .Y(EX__n101) );
  BUFx12f_ASAP7_75t_R EX___U331 ( .A(EX__n1366), .Y(EX__n102) );
  BUFx12f_ASAP7_75t_R EX___U332 ( .A(EX__n394), .Y(EX__n103) );
  BUFx12f_ASAP7_75t_R EX___U333 ( .A(EX__n143), .Y(EX__n926) );
  BUFx16f_ASAP7_75t_R EX___U334 ( .A(EX__n110), .Y(EX__n106) );
  INVx6_ASAP7_75t_R EX___U335 ( .A(EX__n126), .Y(EX__n125) );
  BUFx16f_ASAP7_75t_R EX___U336 ( .A(EX__n1025), .Y(EX__n107) );
  BUFx12f_ASAP7_75t_R EX___U337 ( .A(EX__n353), .Y(EX__n1025) );
  BUFx2_ASAP7_75t_R EX___U338 ( .A(EX__n1421), .Y(EX__n108) );
  BUFx2_ASAP7_75t_R EX___U339 ( .A(EX__n1420), .Y(EX__n109) );
  BUFx12f_ASAP7_75t_R EX___U340 ( .A(EX__n162), .Y(EX__n970) );
  CKINVDCx20_ASAP7_75t_R EX___U341 ( .A(EX__n118), .Y(EX__n112) );
  BUFx12f_ASAP7_75t_R EX___U342 ( .A(EX__n1021), .Y(EX__n126) );
  CKINVDCx9p33_ASAP7_75t_R EX___U343 ( .A(EX__n127), .Y(EX__n389) );
  BUFx16f_ASAP7_75t_R EX___U344 ( .A(EX__n286), .Y(EX__n113) );
  BUFx12f_ASAP7_75t_R EX___U345 ( .A(EX__n781), .Y(EX__n286) );
  CKINVDCx20_ASAP7_75t_R EX___U346 ( .A(EX__n441), .Y(EX__n1222) );
  CKINVDCx20_ASAP7_75t_R EX___U347 ( .A(EX__n107), .Y(EX__n114) );
  BUFx16f_ASAP7_75t_R EX___U348 ( .A(EX__n1069), .Y(EX__n115) );
  BUFx12f_ASAP7_75t_R EX___U349 ( .A(EX__n155), .Y(EX__n1069) );
  BUFx2_ASAP7_75t_R EX___U350 ( .A(EX__n1424), .Y(EX__n116) );
  BUFx2_ASAP7_75t_R EX___U351 ( .A(EX__n1423), .Y(EX__n117) );
  BUFx16f_ASAP7_75t_R EX___U352 ( .A(EX__n125), .Y(EX__n118) );
  BUFx12f_ASAP7_75t_R EX___U353 ( .A(EX__n79), .Y(EX__n119) );
  BUFx12f_ASAP7_75t_R EX___U354 ( .A(EX__n78), .Y(EX__n120) );
  BUFx12f_ASAP7_75t_R EX___U355 ( .A(EX__n1318), .Y(EX__n121) );
  CKINVDCx20_ASAP7_75t_R EX___U356 ( .A(EX__n115), .Y(EX__n122) );
  BUFx2_ASAP7_75t_R EX___U357 ( .A(EX__n1400), .Y(EX__n123) );
  BUFx2_ASAP7_75t_R EX___U358 ( .A(EX__n1399), .Y(EX__n124) );
  BUFx12f_ASAP7_75t_R EX___U359 ( .A(EX__n183), .Y(EX__n1021) );
  BUFx16f_ASAP7_75t_R EX___U360 ( .A(EX__n802), .Y(EX__n127) );
  BUFx12f_ASAP7_75t_R EX___U361 ( .A(EX__n137), .Y(EX__n802) );
  BUFx3_ASAP7_75t_R EX___U362 ( .A(EX__n129), .Y(EX__n128) );
  BUFx2_ASAP7_75t_R EX___U363 ( .A(input_data_2[12]), .Y(EX__n129) );
  BUFx12f_ASAP7_75t_R EX___U364 ( .A(EX__n350), .Y(EX__n130) );
  CKINVDCx20_ASAP7_75t_R EX___U365 ( .A(EX__n861), .Y(EX__n352) );
  BUFx4f_ASAP7_75t_R EX___U366 ( .A(EX__n128), .Y(EX__n351) );
  BUFx2_ASAP7_75t_R EX___U367 ( .A(EX__n1406), .Y(EX__n131) );
  BUFx2_ASAP7_75t_R EX___U368 ( .A(EX__n1405), .Y(EX__n132) );
  BUFx2_ASAP7_75t_R EX___U369 ( .A(EX__n1427), .Y(EX__n133) );
  BUFx2_ASAP7_75t_R EX___U370 ( .A(EX__n1426), .Y(EX__n134) );
  BUFx3_ASAP7_75t_R EX___U371 ( .A(EX__n136), .Y(EX__n135) );
  BUFx2_ASAP7_75t_R EX___U372 ( .A(input_data_2[11]), .Y(EX__n136) );
  BUFx12f_ASAP7_75t_R EX___U373 ( .A(EX__n387), .Y(EX__n137) );
  BUFx4f_ASAP7_75t_R EX___U374 ( .A(EX__n135), .Y(EX__n388) );
  BUFx16f_ASAP7_75t_R EX___U375 ( .A(EX__n1030), .Y(EX__n141) );
  BUFx12f_ASAP7_75t_R EX___U376 ( .A(EX__n539), .Y(EX__n1030) );
  BUFx16f_ASAP7_75t_R EX___U377 ( .A(EX__n930), .Y(EX__n142) );
  BUFx12f_ASAP7_75t_R EX___U378 ( .A(EX__n197), .Y(EX__n930) );
  BUFx12f_ASAP7_75t_R EX___U379 ( .A(input_A[15]), .Y(EX__n143) );
  BUFx4f_ASAP7_75t_R EX___U380 ( .A(EX__n145), .Y(EX__n144) );
  BUFx3_ASAP7_75t_R EX___U381 ( .A(EX__n108), .Y(EX__n145) );
  BUFx4f_ASAP7_75t_R EX___U382 ( .A(EX__n147), .Y(EX__n146) );
  BUFx3_ASAP7_75t_R EX___U383 ( .A(EX__n109), .Y(EX__n147) );
  BUFx3_ASAP7_75t_R EX___U384 ( .A(EX__n150), .Y(EX__n149) );
  BUFx2_ASAP7_75t_R EX___U385 ( .A(input_data_2[6]), .Y(EX__n150) );
  BUFx4f_ASAP7_75t_R EX___U386 ( .A(EX__n149), .Y(EX__n285) );
  BUFx12f_ASAP7_75t_R EX___U387 ( .A(EX__n284), .Y(EX__n781) );
  CKINVDCx20_ASAP7_75t_R EX___U388 ( .A(EX__n142), .Y(EX__n151) );
  BUFx2_ASAP7_75t_R EX___U389 ( .A(EX__n1439), .Y(EX__n152) );
  BUFx2_ASAP7_75t_R EX___U390 ( .A(EX__n1438), .Y(EX__n153) );
  BUFx16f_ASAP7_75t_R EX___U391 ( .A(EX__n974), .Y(EX__n154) );
  BUFx12f_ASAP7_75t_R EX___U392 ( .A(EX__n211), .Y(EX__n974) );
  BUFx12f_ASAP7_75t_R EX___U393 ( .A(input_A[20]), .Y(EX__n155) );
  BUFx4f_ASAP7_75t_R EX___U394 ( .A(EX__n157), .Y(EX__n156) );
  BUFx3_ASAP7_75t_R EX___U395 ( .A(EX__n131), .Y(EX__n157) );
  BUFx4f_ASAP7_75t_R EX___U396 ( .A(EX__n159), .Y(EX__n158) );
  BUFx3_ASAP7_75t_R EX___U397 ( .A(EX__n132), .Y(EX__n159) );
  CKINVDCx20_ASAP7_75t_R EX___U398 ( .A(EX__n122), .Y(EX__n160) );
  CKINVDCx20_ASAP7_75t_R EX___U399 ( .A(EX__n160), .Y(EX__n161) );
  BUFx12f_ASAP7_75t_R EX___U400 ( .A(input_A[14]), .Y(EX__n162) );
  BUFx4f_ASAP7_75t_R EX___U401 ( .A(EX__n164), .Y(EX__n163) );
  BUFx3_ASAP7_75t_R EX___U402 ( .A(EX__n116), .Y(EX__n164) );
  BUFx4f_ASAP7_75t_R EX___U403 ( .A(EX__n166), .Y(EX__n165) );
  BUFx3_ASAP7_75t_R EX___U404 ( .A(EX__n117), .Y(EX__n166) );
  BUFx3_ASAP7_75t_R EX___U405 ( .A(EX__n168), .Y(EX__n167) );
  BUFx2_ASAP7_75t_R EX___U406 ( .A(input_data_2[29]), .Y(EX__n168) );
  BUFx16f_ASAP7_75t_R EX___U407 ( .A(EX__n508), .Y(EX__n169) );
  CKINVDCx10_ASAP7_75t_R EX___U408 ( .A(EX__n169), .Y(EX__n1123) );
  BUFx12f_ASAP7_75t_R EX___U409 ( .A(EX__n509), .Y(EX__n508) );
  CKINVDCx20_ASAP7_75t_R EX___U410 ( .A(EX__n154), .Y(EX__n170) );
  BUFx16f_ASAP7_75t_R EX___U411 ( .A(EX__n1061), .Y(EX__n171) );
  BUFx12f_ASAP7_75t_R EX___U412 ( .A(EX__n235), .Y(EX__n1061) );
  BUFx16f_ASAP7_75t_R EX___U413 ( .A(EX__n921), .Y(EX__n172) );
  BUFx12f_ASAP7_75t_R EX___U414 ( .A(EX__n246), .Y(EX__n921) );
  BUFx2_ASAP7_75t_R EX___U415 ( .A(EX__n1442), .Y(EX__n173) );
  BUFx2_ASAP7_75t_R EX___U416 ( .A(EX__n1441), .Y(EX__n174) );
  BUFx12f_ASAP7_75t_R EX___U417 ( .A(EX__n453), .Y(EX__n175) );
  BUFx3_ASAP7_75t_R EX___U418 ( .A(EX__n177), .Y(EX__n176) );
  BUFx2_ASAP7_75t_R EX___U419 ( .A(input_data_2[28]), .Y(EX__n177) );
  BUFx16f_ASAP7_75t_R EX___U420 ( .A(EX__n477), .Y(EX__n178) );
  INVx13_ASAP7_75t_R EX___U421 ( .A(EX__n178), .Y(EX__n1033) );
  BUFx12f_ASAP7_75t_R EX___U422 ( .A(EX__n478), .Y(EX__n477) );
  CKINVDCx20_ASAP7_75t_R EX___U423 ( .A(EX__n171), .Y(EX__n179) );
  CKINVDCx20_ASAP7_75t_R EX___U424 ( .A(EX__n172), .Y(EX__n180) );
  BUFx2_ASAP7_75t_R EX___U425 ( .A(EX__n1448), .Y(EX__n181) );
  BUFx2_ASAP7_75t_R EX___U426 ( .A(EX__n1447), .Y(EX__n182) );
  BUFx12f_ASAP7_75t_R EX___U427 ( .A(input_A[13]), .Y(EX__n183) );
  BUFx4f_ASAP7_75t_R EX___U428 ( .A(EX__n185), .Y(EX__n184) );
  BUFx3_ASAP7_75t_R EX___U429 ( .A(EX__n133), .Y(EX__n185) );
  BUFx4f_ASAP7_75t_R EX___U430 ( .A(EX__n187), .Y(EX__n186) );
  BUFx3_ASAP7_75t_R EX___U431 ( .A(EX__n134), .Y(EX__n187) );
  BUFx16f_ASAP7_75t_R EX___U432 ( .A(EX__n206), .Y(EX__n188) );
  BUFx12f_ASAP7_75t_R EX___U433 ( .A(EX__n550), .Y(EX__n206) );
  BUFx12f_ASAP7_75t_R EX___U434 ( .A(EX__n175), .Y(EX__n189) );
  BUFx3_ASAP7_75t_R EX___U435 ( .A(EX__n191), .Y(EX__n190) );
  BUFx2_ASAP7_75t_R EX___U436 ( .A(input_data_2[26]), .Y(EX__n191) );
  BUFx2_ASAP7_75t_R EX___U437 ( .A(EX__n1457), .Y(EX__n192) );
  BUFx2_ASAP7_75t_R EX___U438 ( .A(EX__n1456), .Y(EX__n193) );
  BUFx2_ASAP7_75t_R EX___U439 ( .A(EX__n1382), .Y(EX__n194) );
  BUFx2_ASAP7_75t_R EX___U440 ( .A(EX__n1381), .Y(EX__n195) );
  BUFx16f_ASAP7_75t_R EX___U441 ( .A(EX__n1161), .Y(EX__n196) );
  BUFx12f_ASAP7_75t_R EX___U442 ( .A(EX__n277), .Y(EX__n1161) );
  BUFx12f_ASAP7_75t_R EX___U443 ( .A(input_A[8]), .Y(EX__n197) );
  BUFx4f_ASAP7_75t_R EX___U444 ( .A(EX__n199), .Y(EX__n198) );
  BUFx3_ASAP7_75t_R EX___U445 ( .A(EX__n173), .Y(EX__n199) );
  BUFx4f_ASAP7_75t_R EX___U446 ( .A(EX__n201), .Y(EX__n200) );
  BUFx3_ASAP7_75t_R EX___U447 ( .A(EX__n174), .Y(EX__n201) );
  CKINVDCx20_ASAP7_75t_R EX___U448 ( .A(EX__n151), .Y(EX__n202) );
  CKINVDCx20_ASAP7_75t_R EX___U449 ( .A(EX__n202), .Y(EX__n203) );
  CKINVDCx9p33_ASAP7_75t_R EX___U450 ( .A(EX__n227), .Y(EX__n341) );
  BUFx3_ASAP7_75t_R EX___U451 ( .A(EX__n205), .Y(EX__n204) );
  BUFx2_ASAP7_75t_R EX___U452 ( .A(input_data_2[10]), .Y(EX__n205) );
  BUFx12f_ASAP7_75t_R EX___U453 ( .A(EX__n551), .Y(EX__n550) );
  CKINVDCx20_ASAP7_75t_R EX___U454 ( .A(EX__n196), .Y(EX__n207) );
  CKINVDCx20_ASAP7_75t_R EX___U455 ( .A(EX__n210), .Y(EX__n208) );
  CKINVDCx20_ASAP7_75t_R EX___U456 ( .A(EX__n208), .Y(EX__n209) );
  BUFx16f_ASAP7_75t_R EX___U457 ( .A(EX__n1016), .Y(EX__n210) );
  BUFx12f_ASAP7_75t_R EX___U458 ( .A(EX__n371), .Y(EX__n1016) );
  BUFx12f_ASAP7_75t_R EX___U459 ( .A(input_A[6]), .Y(EX__n211) );
  BUFx4f_ASAP7_75t_R EX___U460 ( .A(EX__n213), .Y(EX__n212) );
  BUFx3_ASAP7_75t_R EX___U461 ( .A(EX__n181), .Y(EX__n213) );
  BUFx4f_ASAP7_75t_R EX___U462 ( .A(EX__n215), .Y(EX__n214) );
  BUFx3_ASAP7_75t_R EX___U463 ( .A(EX__n182), .Y(EX__n215) );
  CKINVDCx20_ASAP7_75t_R EX___U464 ( .A(EX__n170), .Y(EX__n216) );
  CKINVDCx20_ASAP7_75t_R EX___U465 ( .A(EX__n216), .Y(EX__n217) );
  CKINVDCx14_ASAP7_75t_R EX___U466 ( .A(EX__n242), .Y(EX__n435) );
  BUFx3_ASAP7_75t_R EX___U467 ( .A(EX__n219), .Y(EX__n218) );
  BUFx2_ASAP7_75t_R EX___U468 ( .A(input_data_2[9]), .Y(EX__n219) );
  BUFx16f_ASAP7_75t_R EX___U469 ( .A(EX__n526), .Y(EX__n220) );
  CKINVDCx10_ASAP7_75t_R EX___U470 ( .A(EX__n220), .Y(EX__n1208) );
  BUFx12f_ASAP7_75t_R EX___U471 ( .A(EX__n527), .Y(EX__n526) );
  BUFx2_ASAP7_75t_R EX___U472 ( .A(EX__n1463), .Y(EX__n221) );
  BUFx2_ASAP7_75t_R EX___U473 ( .A(EX__n1462), .Y(EX__n222) );
  BUFx2_ASAP7_75t_R EX___U474 ( .A(EX__n1385), .Y(EX__n223) );
  BUFx2_ASAP7_75t_R EX___U475 ( .A(EX__n1384), .Y(EX__n224) );
  CKINVDCx20_ASAP7_75t_R EX___U476 ( .A(EX__n226), .Y(EX__n225) );
  BUFx16f_ASAP7_75t_R EX___U477 ( .A(EX__n1110), .Y(EX__n226) );
  BUFx16f_ASAP7_75t_R EX___U478 ( .A(EX__n821), .Y(EX__n227) );
  BUFx12f_ASAP7_75t_R EX___U479 ( .A(EX__n245), .Y(EX__n821) );
  BUFx3_ASAP7_75t_R EX___U480 ( .A(EX__n229), .Y(EX__n228) );
  BUFx2_ASAP7_75t_R EX___U481 ( .A(input_data_2[8]), .Y(EX__n229) );
  BUFx12f_ASAP7_75t_R EX___U482 ( .A(EX__n617), .Y(EX__n230) );
  BUFx2_ASAP7_75t_R EX___U483 ( .A(EX__n1430), .Y(EX__n231) );
  BUFx2_ASAP7_75t_R EX___U484 ( .A(EX__n1429), .Y(EX__n232) );
  CKINVDCx20_ASAP7_75t_R EX___U485 ( .A(EX__n225), .Y(EX__n233) );
  CKINVDCx20_ASAP7_75t_R EX___U486 ( .A(EX__n233), .Y(EX__n234) );
  BUFx12f_ASAP7_75t_R EX___U487 ( .A(EX__n299), .Y(EX__n1110) );
  BUFx12f_ASAP7_75t_R EX___U488 ( .A(input_A[3]), .Y(EX__n235) );
  BUFx4f_ASAP7_75t_R EX___U489 ( .A(EX__n237), .Y(EX__n236) );
  BUFx3_ASAP7_75t_R EX___U490 ( .A(EX__n192), .Y(EX__n237) );
  BUFx4f_ASAP7_75t_R EX___U491 ( .A(EX__n239), .Y(EX__n238) );
  BUFx3_ASAP7_75t_R EX___U492 ( .A(EX__n193), .Y(EX__n239) );
  CKINVDCx20_ASAP7_75t_R EX___U493 ( .A(EX__n179), .Y(EX__n240) );
  CKINVDCx20_ASAP7_75t_R EX___U494 ( .A(EX__n240), .Y(EX__n241) );
  BUFx16f_ASAP7_75t_R EX___U495 ( .A(EX__n260), .Y(EX__n242) );
  BUFx12f_ASAP7_75t_R EX___U496 ( .A(EX__n261), .Y(EX__n260) );
  BUFx3_ASAP7_75t_R EX___U497 ( .A(EX__n244), .Y(EX__n243) );
  BUFx2_ASAP7_75t_R EX___U498 ( .A(input_data_2[7]), .Y(EX__n244) );
  BUFx12f_ASAP7_75t_R EX___U499 ( .A(EX__n339), .Y(EX__n245) );
  BUFx4f_ASAP7_75t_R EX___U500 ( .A(EX__n243), .Y(EX__n340) );
  INVx6_ASAP7_75t_R EX___U501 ( .A(EX__n276), .Y(EX__n275) );
  BUFx12f_ASAP7_75t_R EX___U502 ( .A(input_A[28]), .Y(EX__n246) );
  BUFx4f_ASAP7_75t_R EX___U503 ( .A(EX__n248), .Y(EX__n247) );
  BUFx3_ASAP7_75t_R EX___U504 ( .A(EX__n194), .Y(EX__n248) );
  BUFx4f_ASAP7_75t_R EX___U505 ( .A(EX__n250), .Y(EX__n249) );
  BUFx3_ASAP7_75t_R EX___U506 ( .A(EX__n195), .Y(EX__n250) );
  CKINVDCx20_ASAP7_75t_R EX___U507 ( .A(EX__n180), .Y(EX__n251) );
  CKINVDCx20_ASAP7_75t_R EX___U508 ( .A(EX__n251), .Y(EX__n252) );
  BUFx12f_ASAP7_75t_R EX___U509 ( .A(EX__n100), .Y(EX__n1364) );
  BUFx12f_ASAP7_75t_R EX___U510 ( .A(EX__n83), .Y(EX__n1358) );
  BUFx12f_ASAP7_75t_R EX___U511 ( .A(EX__n290), .Y(EX__n253) );
  BUFx2_ASAP7_75t_R EX___U512 ( .A(EX__n1349), .Y(EX__n254) );
  BUFx12f_ASAP7_75t_R EX___U513 ( .A(EX__n1349), .Y(EX__n255) );
  BUFx2_ASAP7_75t_R EX___U514 ( .A(EX__n1349), .Y(EX__n256) );
  BUFx2_ASAP7_75t_R EX___U515 ( .A(EX__n1349), .Y(EX__n257) );
  BUFx16f_ASAP7_75t_R EX___U516 ( .A(EX__n1065), .Y(EX__n258) );
  BUFx12f_ASAP7_75t_R EX___U517 ( .A(EX__n376), .Y(EX__n1065) );
  CKINVDCx20_ASAP7_75t_R EX___U518 ( .A(EX__n271), .Y(EX__n259) );
  BUFx12f_ASAP7_75t_R EX___U519 ( .A(EX__n1074), .Y(EX__n276) );
  BUFx12f_ASAP7_75t_R EX___U520 ( .A(EX__n272), .Y(EX__n261) );
  BUFx10_ASAP7_75t_R EX___U521 ( .A(input_data_2[27]), .Y(EX__n272) );
  BUFx2_ASAP7_75t_R EX___U522 ( .A(EX__n1344), .Y(EX__n262) );
  BUFx12f_ASAP7_75t_R EX___U523 ( .A(EX__n1344), .Y(EX__n263) );
  BUFx2_ASAP7_75t_R EX___U524 ( .A(EX__n1344), .Y(EX__n264) );
  BUFx2_ASAP7_75t_R EX___U525 ( .A(EX__n1344), .Y(EX__n265) );
  BUFx12f_ASAP7_75t_R EX___U526 ( .A(EX__n287), .Y(EX__n266) );
  BUFx12f_ASAP7_75t_R EX___U527 ( .A(EX__n287), .Y(EX__n267) );
  BUFx12f_ASAP7_75t_R EX___U528 ( .A(EX__n269), .Y(EX__n268) );
  BUFx12f_ASAP7_75t_R EX___U529 ( .A(EX__n402), .Y(EX__n269) );
  BUFx12f_ASAP7_75t_R EX___U530 ( .A(EX__n291), .Y(EX__n270) );
  BUFx16f_ASAP7_75t_R EX___U531 ( .A(EX__n275), .Y(EX__n271) );
  BUFx12f_ASAP7_75t_R EX___U532 ( .A(EX__n295), .Y(EX__n273) );
  CKINVDCx20_ASAP7_75t_R EX___U533 ( .A(EX__n258), .Y(EX__n274) );
  BUFx12f_ASAP7_75t_R EX___U534 ( .A(EX__n326), .Y(EX__n1074) );
  BUFx12f_ASAP7_75t_R EX___U535 ( .A(input_A[27]), .Y(EX__n277) );
  BUFx4f_ASAP7_75t_R EX___U536 ( .A(EX__n279), .Y(EX__n278) );
  BUFx3_ASAP7_75t_R EX___U537 ( .A(EX__n223), .Y(EX__n279) );
  BUFx4f_ASAP7_75t_R EX___U538 ( .A(EX__n281), .Y(EX__n280) );
  BUFx3_ASAP7_75t_R EX___U539 ( .A(EX__n224), .Y(EX__n281) );
  CKINVDCx20_ASAP7_75t_R EX___U540 ( .A(EX__n207), .Y(EX__n282) );
  CKINVDCx20_ASAP7_75t_R EX___U541 ( .A(EX__n282), .Y(EX__n283) );
  BUFx6f_ASAP7_75t_R EX___U542 ( .A(EX__n285), .Y(EX__n284) );
  BUFx12f_ASAP7_75t_R EX___U543 ( .A(EX__n1368), .Y(EX__n287) );
  BUFx12f_ASAP7_75t_R EX___U544 ( .A(EX__n403), .Y(EX__n288) );
  BUFx12f_ASAP7_75t_R EX___U545 ( .A(EX__n288), .Y(EX__n289) );
  BUFx12f_ASAP7_75t_R EX___U546 ( .A(EX__n1341), .Y(EX__n290) );
  BUFx12f_ASAP7_75t_R EX___U547 ( .A(EX__n325), .Y(EX__n291) );
  BUFx16f_ASAP7_75t_R EX___U548 ( .A(EX__n965), .Y(EX__n292) );
  BUFx12f_ASAP7_75t_R EX___U549 ( .A(EX__n446), .Y(EX__n965) );
  BUFx3_ASAP7_75t_R EX___U550 ( .A(EX__n294), .Y(EX__n293) );
  BUFx2_ASAP7_75t_R EX___U551 ( .A(EX__n1469), .Y(EX__n294) );
  BUFx12f_ASAP7_75t_R EX___U552 ( .A(EX__n314), .Y(EX__n295) );
  BUFx2_ASAP7_75t_R EX___U553 ( .A(EX__n1466), .Y(EX__n296) );
  BUFx2_ASAP7_75t_R EX___U554 ( .A(EX__n1465), .Y(EX__n297) );
  BUFx16f_ASAP7_75t_R EX___U555 ( .A(EX__n1101), .Y(EX__n298) );
  BUFx12f_ASAP7_75t_R EX___U556 ( .A(EX__n495), .Y(EX__n1101) );
  CKINVDCx14_ASAP7_75t_R EX___U557 ( .A(EX__n490), .Y(EX__n1162) );
  CKINVDCx14_ASAP7_75t_R EX___U558 ( .A(EX__n1077), .Y(EX__n619) );
  BUFx12f_ASAP7_75t_R EX___U559 ( .A(input_A[12]), .Y(EX__n299) );
  BUFx4f_ASAP7_75t_R EX___U560 ( .A(EX__n301), .Y(EX__n300) );
  BUFx3_ASAP7_75t_R EX___U561 ( .A(EX__n231), .Y(EX__n301) );
  BUFx4f_ASAP7_75t_R EX___U562 ( .A(EX__n303), .Y(EX__n302) );
  BUFx3_ASAP7_75t_R EX___U563 ( .A(EX__n232), .Y(EX__n303) );
  CKINVDCx20_ASAP7_75t_R EX___U564 ( .A(EX__n305), .Y(EX__n304) );
  BUFx16f_ASAP7_75t_R EX___U565 ( .A(EX__n1226), .Y(EX__n305) );
  BUFx12f_ASAP7_75t_R EX___U566 ( .A(EX__n313), .Y(EX__n306) );
  BUFx12f_ASAP7_75t_R EX___U567 ( .A(EX__n313), .Y(EX__n307) );
  CKINVDCx14_ASAP7_75t_R EX___U568 ( .A(EX__n1219), .Y(EX__n858) );
  BUFx12f_ASAP7_75t_R EX___U569 ( .A(EX__n310), .Y(EX__n308) );
  BUFx12f_ASAP7_75t_R EX___U570 ( .A(EX__n311), .Y(EX__n309) );
  BUFx12f_ASAP7_75t_R EX___U571 ( .A(EX__n80), .Y(EX__n310) );
  BUFx12f_ASAP7_75t_R EX___U572 ( .A(EX__n80), .Y(EX__n311) );
  BUFx6f_ASAP7_75t_R EX___U573 ( .A(EX__n309), .Y(EX__n1300) );
  BUFx12f_ASAP7_75t_R EX___U574 ( .A(EX__n1306), .Y(EX__n1304) );
  BUFx16f_ASAP7_75t_R EX___U575 ( .A(EX__n322), .Y(EX__n312) );
  BUFx12f_ASAP7_75t_R EX___U576 ( .A(EX__n398), .Y(EX__n322) );
  BUFx12f_ASAP7_75t_R EX___U577 ( .A(EX__n331), .Y(EX__n1226) );
  BUFx12f_ASAP7_75t_R EX___U578 ( .A(EX__n437), .Y(EX__n313) );
  BUFx12f_ASAP7_75t_R EX___U579 ( .A(EX__n1263), .Y(EX__n314) );
  CKINVDCx20_ASAP7_75t_R EX___U580 ( .A(EX__n298), .Y(EX__n315) );
  BUFx2_ASAP7_75t_R EX___U581 ( .A(EX__n1394), .Y(EX__n316) );
  BUFx2_ASAP7_75t_R EX___U582 ( .A(EX__n1393), .Y(EX__n317) );
  BUFx2_ASAP7_75t_R EX___U583 ( .A(EX__n1418), .Y(EX__n318) );
  BUFx2_ASAP7_75t_R EX___U584 ( .A(EX__n1417), .Y(EX__n319) );
  BUFx6f_ASAP7_75t_R EX___U585 ( .A(EX__n1302), .Y(EX__n1297) );
  BUFx6f_ASAP7_75t_R EX___U586 ( .A(EX__n362), .Y(EX__n1296) );
  BUFx6f_ASAP7_75t_R EX___U587 ( .A(EX__n1303), .Y(EX__n1295) );
  CKINVDCx20_ASAP7_75t_R EX___U588 ( .A(EX__n312), .Y(EX__n320) );
  CKINVDCx20_ASAP7_75t_R EX___U589 ( .A(EX__n320), .Y(EX__n321) );
  INVx5_ASAP7_75t_R EX___U590 ( .A(EX__n1234), .Y(EX__n398) );
  BUFx12f_ASAP7_75t_R EX___U591 ( .A(EX__n607), .Y(EX__n323) );
  BUFx12f_ASAP7_75t_R EX___U592 ( .A(EX__n607), .Y(EX__n324) );
  BUFx12f_ASAP7_75t_R EX___U593 ( .A(EX__n457), .Y(EX__n325) );
  CKINVDCx14_ASAP7_75t_R EX___U594 ( .A(EX__n1031), .Y(EX__n701) );
  BUFx12f_ASAP7_75t_R EX___U595 ( .A(input_A[16]), .Y(EX__n326) );
  BUFx4f_ASAP7_75t_R EX___U596 ( .A(EX__n328), .Y(EX__n327) );
  BUFx3_ASAP7_75t_R EX___U597 ( .A(EX__n318), .Y(EX__n328) );
  BUFx4f_ASAP7_75t_R EX___U598 ( .A(EX__n330), .Y(EX__n329) );
  BUFx3_ASAP7_75t_R EX___U599 ( .A(EX__n319), .Y(EX__n330) );
  BUFx12f_ASAP7_75t_R EX___U600 ( .A(input_A[21]), .Y(EX__n331) );
  CKINVDCx20_ASAP7_75t_R EX___U601 ( .A(EX__n304), .Y(EX__n332) );
  CKINVDCx20_ASAP7_75t_R EX___U602 ( .A(EX__n332), .Y(EX__n333) );
  BUFx2_ASAP7_75t_R EX___U603 ( .A(EX__n1403), .Y(EX__n334) );
  BUFx2_ASAP7_75t_R EX___U604 ( .A(EX__n1402), .Y(EX__n335) );
  CKINVDCx20_ASAP7_75t_R EX___U605 ( .A(EX__n337), .Y(EX__n336) );
  BUFx16f_ASAP7_75t_R EX___U606 ( .A(EX__n1183), .Y(EX__n337) );
  BUFx16f_ASAP7_75t_R EX___U607 ( .A(EX__n349), .Y(EX__n338) );
  BUFx12f_ASAP7_75t_R EX___U608 ( .A(EX__n384), .Y(EX__n349) );
  BUFx6f_ASAP7_75t_R EX___U609 ( .A(EX__n340), .Y(EX__n339) );
  BUFx12f_ASAP7_75t_R EX___U610 ( .A(EX__n456), .Y(EX__n342) );
  BUFx12f_ASAP7_75t_R EX___U611 ( .A(EX__n456), .Y(EX__n343) );
  BUFx12f_ASAP7_75t_R EX___U612 ( .A(EX__n480), .Y(EX__n344) );
  BUFx2_ASAP7_75t_R EX___U613 ( .A(EX__n1388), .Y(EX__n345) );
  BUFx2_ASAP7_75t_R EX___U614 ( .A(EX__n1387), .Y(EX__n346) );
  BUFx12f_ASAP7_75t_R EX___U615 ( .A(EX__n364), .Y(EX__n1183) );
  CKINVDCx20_ASAP7_75t_R EX___U616 ( .A(EX__n338), .Y(EX__n347) );
  CKINVDCx20_ASAP7_75t_R EX___U617 ( .A(EX__n347), .Y(EX__n348) );
  INVx5_ASAP7_75t_R EX___U618 ( .A(EX__n1230), .Y(EX__n384) );
  BUFx6f_ASAP7_75t_R EX___U619 ( .A(EX__n351), .Y(EX__n350) );
  BUFx16f_ASAP7_75t_R EX___U620 ( .A(EX__n130), .Y(EX__n861) );
  BUFx12f_ASAP7_75t_R EX___U621 ( .A(input_A[22]), .Y(EX__n353) );
  BUFx4f_ASAP7_75t_R EX___U622 ( .A(EX__n355), .Y(EX__n354) );
  BUFx3_ASAP7_75t_R EX___U623 ( .A(EX__n123), .Y(EX__n355) );
  BUFx4f_ASAP7_75t_R EX___U624 ( .A(EX__n357), .Y(EX__n356) );
  BUFx3_ASAP7_75t_R EX___U625 ( .A(EX__n124), .Y(EX__n357) );
  CKINVDCx20_ASAP7_75t_R EX___U626 ( .A(EX__n114), .Y(EX__n358) );
  CKINVDCx20_ASAP7_75t_R EX___U627 ( .A(EX__n358), .Y(EX__n359) );
  BUFx12f_ASAP7_75t_R EX___U628 ( .A(EX__n362), .Y(EX__n360) );
  BUFx12f_ASAP7_75t_R EX___U629 ( .A(EX__n363), .Y(EX__n361) );
  BUFx12f_ASAP7_75t_R EX___U630 ( .A(EX__n1305), .Y(EX__n362) );
  BUFx12f_ASAP7_75t_R EX___U631 ( .A(EX__n1308), .Y(EX__n363) );
  BUFx12f_ASAP7_75t_R EX___U632 ( .A(EX__n1301), .Y(EX__n1308) );
  BUFx12f_ASAP7_75t_R EX___U633 ( .A(input_A[18]), .Y(EX__n364) );
  CKINVDCx20_ASAP7_75t_R EX___U634 ( .A(EX__n336), .Y(EX__n365) );
  CKINVDCx20_ASAP7_75t_R EX___U635 ( .A(EX__n365), .Y(EX__n366) );
  BUFx2_ASAP7_75t_R EX___U636 ( .A(EX__n1412), .Y(EX__n367) );
  BUFx2_ASAP7_75t_R EX___U637 ( .A(EX__n1411), .Y(EX__n368) );
  CKINVDCx10_ASAP7_75t_R EX___U638 ( .A(EX__n461), .Y(EX__n777) );
  INVx6_ASAP7_75t_R EX___U639 ( .A(EX__n420), .Y(EX__n408) );
  BUFx16f_ASAP7_75t_R EX___U640 ( .A(EX__n1011), .Y(EX__n370) );
  BUFx12f_ASAP7_75t_R EX___U641 ( .A(EX__n593), .Y(EX__n1011) );
  BUFx12f_ASAP7_75t_R EX___U642 ( .A(input_A[1]), .Y(EX__n371) );
  BUFx4f_ASAP7_75t_R EX___U643 ( .A(EX__n373), .Y(EX__n372) );
  BUFx3_ASAP7_75t_R EX___U644 ( .A(EX__n221), .Y(EX__n373) );
  BUFx4f_ASAP7_75t_R EX___U645 ( .A(EX__n375), .Y(EX__n374) );
  BUFx3_ASAP7_75t_R EX___U646 ( .A(EX__n222), .Y(EX__n375) );
  BUFx12f_ASAP7_75t_R EX___U647 ( .A(input_A[24]), .Y(EX__n376) );
  BUFx4f_ASAP7_75t_R EX___U648 ( .A(EX__n378), .Y(EX__n377) );
  BUFx3_ASAP7_75t_R EX___U649 ( .A(EX__n316), .Y(EX__n378) );
  BUFx4f_ASAP7_75t_R EX___U650 ( .A(EX__n380), .Y(EX__n379) );
  BUFx3_ASAP7_75t_R EX___U651 ( .A(EX__n317), .Y(EX__n380) );
  CKINVDCx20_ASAP7_75t_R EX___U652 ( .A(EX__n274), .Y(EX__n381) );
  CKINVDCx20_ASAP7_75t_R EX___U653 ( .A(EX__n381), .Y(EX__n382) );
  BUFx12f_ASAP7_75t_R EX___U654 ( .A(input_A[10]), .Y(EX__n383) );
  BUFx2_ASAP7_75t_R EX___U655 ( .A(EX__n1436), .Y(EX__n385) );
  BUFx2_ASAP7_75t_R EX___U656 ( .A(EX__n1435), .Y(EX__n386) );
  BUFx6f_ASAP7_75t_R EX___U657 ( .A(EX__n388), .Y(EX__n387) );
  BUFx16f_ASAP7_75t_R EX___U658 ( .A(EX__n408), .Y(EX__n391) );
  BUFx12f_ASAP7_75t_R EX___U659 ( .A(EX__n1092), .Y(EX__n420) );
  BUFx2_ASAP7_75t_R EX___U660 ( .A(EX__n1376), .Y(EX__n392) );
  BUFx2_ASAP7_75t_R EX___U661 ( .A(EX__n1375), .Y(EX__n393) );
  BUFx12f_ASAP7_75t_R EX___U662 ( .A(EX__n1320), .Y(EX__n394) );
  BUFx12f_ASAP7_75t_R EX___U663 ( .A(EX__n396), .Y(EX__n395) );
  INVx4_ASAP7_75t_R EX___U664 ( .A(EX__n360), .Y(EX__n396) );
  BUFx12f_ASAP7_75t_R EX___U665 ( .A(ID_EX_ALUSrc), .Y(EX__n1320) );
  BUFx12f_ASAP7_75t_R EX___U666 ( .A(input_A[5]), .Y(EX__n397) );
  BUFx2_ASAP7_75t_R EX___U667 ( .A(EX__n1451), .Y(EX__n399) );
  BUFx2_ASAP7_75t_R EX___U668 ( .A(EX__n1450), .Y(EX__n400) );
  BUFx12f_ASAP7_75t_R EX___U669 ( .A(EX__n1369), .Y(EX__n401) );
  BUFx12f_ASAP7_75t_R EX___U670 ( .A(EX__n460), .Y(EX__n402) );
  BUFx12f_ASAP7_75t_R EX___U671 ( .A(EX__n514), .Y(EX__n403) );
  BUFx12f_ASAP7_75t_R EX___U672 ( .A(EX__n95), .Y(EX__n406) );
  BUFx12f_ASAP7_75t_R EX___U673 ( .A(EX__n94), .Y(EX__n407) );
  BUFx12f_ASAP7_75t_R EX___U674 ( .A(EX__n395), .Y(EX__n1317) );
  BUFx12f_ASAP7_75t_R EX___U675 ( .A(EX__n77), .Y(EX__n1318) );
  BUFx12f_ASAP7_75t_R EX___U676 ( .A(EX__n76), .Y(EX__n1319) );
  CKINVDCx12_ASAP7_75t_R EX___U677 ( .A(EX__n427), .Y(EX__n637) );
  INVx6_ASAP7_75t_R EX___U678 ( .A(EX__n463), .Y(EX__n462) );
  CKINVDCx20_ASAP7_75t_R EX___U679 ( .A(EX__n391), .Y(EX__n409) );
  CKINVDCx16_ASAP7_75t_R EX___U680 ( .A(EX__n1170), .Y(EX__n794) );
  BUFx6f_ASAP7_75t_R EX___U681 ( .A(EX__n1316), .Y(EX__n1315) );
  BUFx6f_ASAP7_75t_R EX___U682 ( .A(EX__n1316), .Y(EX__n1314) );
  BUFx12f_ASAP7_75t_R EX___U683 ( .A(EX__n1321), .Y(EX__n1316) );
  CKINVDCx9p33_ASAP7_75t_R EX___U684 ( .A(EX__n468), .Y(EX__n960) );
  INVx6_ASAP7_75t_R EX___U685 ( .A(EX__n471), .Y(EX__n469) );
  BUFx3_ASAP7_75t_R EX___U686 ( .A(EX__n369), .Y(EX__n415) );
  BUFx3_ASAP7_75t_R EX___U687 ( .A(EX__n417), .Y(EX__n416) );
  BUFx2_ASAP7_75t_R EX___U688 ( .A(EX__n1562), .Y(EX__n417) );
  BUFx2_ASAP7_75t_R EX___U689 ( .A(EX__n1373), .Y(EX__n418) );
  BUFx2_ASAP7_75t_R EX___U690 ( .A(EX__n1372), .Y(EX__n419) );
  BUFx12f_ASAP7_75t_R EX___U691 ( .A(EX__n503), .Y(EX__n1092) );
  BUFx16f_ASAP7_75t_R EX___U692 ( .A(EX__n451), .Y(EX__n421) );
  INVx13_ASAP7_75t_R EX___U693 ( .A(EX__n421), .Y(EX__n427) );
  BUFx12f_ASAP7_75t_R EX___U694 ( .A(EX__n502), .Y(EX__n451) );
  BUFx12f_ASAP7_75t_R EX___U695 ( .A(ALU_ctl[2]), .Y(EX__n422) );
  BUFx12f_ASAP7_75t_R EX___U696 ( .A(EX__n1307), .Y(EX__n1305) );
  BUFx12f_ASAP7_75t_R EX___U697 ( .A(EX__n1307), .Y(EX__n1306) );
  BUFx12f_ASAP7_75t_R EX___U698 ( .A(EX__n361), .Y(EX__n1307) );
  BUFx3_ASAP7_75t_R EX___U699 ( .A(EX__n1036), .Y(EX__n1035) );
  BUFx12f_ASAP7_75t_R EX___U700 ( .A(EX__n808), .Y(EX__n423) );
  BUFx3_ASAP7_75t_R EX___U701 ( .A(EX__n425), .Y(EX__n424) );
  BUFx2_ASAP7_75t_R EX___U702 ( .A(input_data_2[18]), .Y(EX__n425) );
  BUFx12f_ASAP7_75t_R EX___U703 ( .A(EX__n856), .Y(EX__n426) );
  BUFx16f_ASAP7_75t_R EX___U704 ( .A(EX__n1175), .Y(EX__n428) );
  BUFx12f_ASAP7_75t_R EX___U705 ( .A(EX__n598), .Y(EX__n1175) );
  BUFx12f_ASAP7_75t_R EX___U706 ( .A(input_A[29]), .Y(EX__n429) );
  CKINVDCx20_ASAP7_75t_R EX___U707 ( .A(EX__n1214), .Y(EX__n430) );
  CKINVDCx20_ASAP7_75t_R EX___U708 ( .A(EX__n430), .Y(EX__n431) );
  BUFx2_ASAP7_75t_R EX___U709 ( .A(EX__n1379), .Y(EX__n432) );
  BUFx2_ASAP7_75t_R EX___U710 ( .A(EX__n1378), .Y(EX__n433) );
  BUFx2_ASAP7_75t_R EX___U711 ( .A(EX__n669), .Y(EX__n436) );
  INVx13_ASAP7_75t_R EX___U712 ( .A(EX__n1237), .Y(EX__n1238) );
  CKINVDCx16_ASAP7_75t_R EX___U713 ( .A(EX__n1211), .Y(EX__n955) );
  BUFx12f_ASAP7_75t_R EX___U714 ( .A(EX__n1279), .Y(EX__n437) );
  BUFx2_ASAP7_75t_R EX___U715 ( .A(EX__n1575), .Y(EX__n438) );
  BUFx3_ASAP7_75t_R EX___U716 ( .A(EX__n440), .Y(EX__n439) );
  BUFx2_ASAP7_75t_R EX___U717 ( .A(input_data_2[15]), .Y(EX__n440) );
  BUFx16f_ASAP7_75t_R EX___U718 ( .A(EX__n809), .Y(EX__n441) );
  BUFx12f_ASAP7_75t_R EX___U719 ( .A(EX__n810), .Y(EX__n809) );
  BUFx16f_ASAP7_75t_R EX___U720 ( .A(EX__n1118), .Y(EX__n442) );
  BUFx12f_ASAP7_75t_R EX___U721 ( .A(EX__n538), .Y(EX__n1118) );
  BUFx3_ASAP7_75t_R EX___U722 ( .A(EX__n444), .Y(EX__n443) );
  BUFx2_ASAP7_75t_R EX___U723 ( .A(input_data_2[17]), .Y(EX__n444) );
  BUFx12f_ASAP7_75t_R EX___U724 ( .A(EX__n788), .Y(EX__n445) );
  BUFx12f_ASAP7_75t_R EX___U725 ( .A(input_A[0]), .Y(EX__n446) );
  BUFx4f_ASAP7_75t_R EX___U726 ( .A(EX__n448), .Y(EX__n447) );
  BUFx3_ASAP7_75t_R EX___U727 ( .A(EX__n296), .Y(EX__n448) );
  BUFx4f_ASAP7_75t_R EX___U728 ( .A(EX__n450), .Y(EX__n449) );
  BUFx3_ASAP7_75t_R EX___U729 ( .A(EX__n297), .Y(EX__n450) );
  BUFx16f_ASAP7_75t_R EX___U730 ( .A(EX__n1186), .Y(EX__n502) );
  CKINVDCx16_ASAP7_75t_R EX___U731 ( .A(EX__n1249), .Y(EX__n552) );
  INVx13_ASAP7_75t_R EX___U732 ( .A(EX__n552), .Y(EX__n553) );
  BUFx16f_ASAP7_75t_R EX___U733 ( .A(EX__n189), .Y(EX__n452) );
  BUFx4f_ASAP7_75t_R EX___U734 ( .A(EX__n190), .Y(EX__n453) );
  BUFx3_ASAP7_75t_R EX___U735 ( .A(EX_read_reg_data_2[26]), .Y(EX__n1490) );
  CKINVDCx10_ASAP7_75t_R EX___U736 ( .A(EX__n452), .Y(EX__n978) );
  BUFx2_ASAP7_75t_R EX___U737 ( .A(EX__n992), .Y(EX__n454) );
  BUFx12f_ASAP7_75t_R EX___U738 ( .A(EX__n343), .Y(EX__n455) );
  BUFx12f_ASAP7_75t_R EX___U739 ( .A(EX__n627), .Y(EX__n456) );
  BUFx12f_ASAP7_75t_R EX___U740 ( .A(EX__n761), .Y(EX__n457) );
  BUFx12f_ASAP7_75t_R EX___U741 ( .A(EX__n459), .Y(EX__n458) );
  BUFx12f_ASAP7_75t_R EX___U742 ( .A(EX__n1353), .Y(EX__n459) );
  BUFx12f_ASAP7_75t_R EX___U743 ( .A(EX__n1338), .Y(EX__n460) );
  BUFx16f_ASAP7_75t_R EX___U744 ( .A(EX__n898), .Y(EX__n461) );
  BUFx12f_ASAP7_75t_R EX___U745 ( .A(EX__n524), .Y(EX__n898) );
  CKINVDCx16_ASAP7_75t_R EX___U746 ( .A(EX__n566), .Y(EX__n798) );
  BUFx12f_ASAP7_75t_R EX___U747 ( .A(EX__n464), .Y(EX__n463) );
  BUFx12f_ASAP7_75t_R EX___U748 ( .A(EX__n138), .Y(EX__n464) );
  AND2x6_ASAP7_75t_R EX___U749 ( .A(EX__n1578), .B(ForwardA[0]), .Y(EX__n138) );
  BUFx3_ASAP7_75t_R EX___U750 ( .A(EX__n466), .Y(EX__n465) );
  BUFx2_ASAP7_75t_R EX___U751 ( .A(input_data_2[30]), .Y(EX__n466) );
  BUFx12f_ASAP7_75t_R EX___U752 ( .A(EX__n957), .Y(EX__n467) );
  BUFx16f_ASAP7_75t_R EX___U753 ( .A(EX__n1167), .Y(EX__n468) );
  BUFx12f_ASAP7_75t_R EX___U754 ( .A(EX__n467), .Y(EX__n1167) );
  BUFx16f_ASAP7_75t_R EX___U755 ( .A(EX__n469), .Y(EX__n546) );
  CKINVDCx14_ASAP7_75t_R EX___U756 ( .A(EX__n546), .Y(EX__n470) );
  BUFx12f_ASAP7_75t_R EX___U757 ( .A(EX__n472), .Y(EX__n471) );
  BUFx12f_ASAP7_75t_R EX___U758 ( .A(EX__n977), .Y(EX__n472) );
  BUFx3_ASAP7_75t_R EX___U759 ( .A(EX__n549), .Y(EX__n473) );
  BUFx6f_ASAP7_75t_R EX___U760 ( .A(EX__n548), .Y(EX__n977) );
  BUFx4f_ASAP7_75t_R EX___U761 ( .A(EX__n473), .Y(EX__n548) );
  BUFx6f_ASAP7_75t_R EX___U762 ( .A(EX__n475), .Y(EX__n474) );
  BUFx4f_ASAP7_75t_R EX___U763 ( .A(EX__n293), .Y(EX__n475) );
  BUFx12f_ASAP7_75t_R EX___U764 ( .A(EX__n474), .Y(EX__n887) );
  INVx5_ASAP7_75t_R EX___U765 ( .A(EX__n887), .Y(EX__n476) );
  AND2x6_ASAP7_75t_R EX___U766 ( .A(EX__n1288), .B(EX__n1572), .Y(EX__n808) );
  BUFx12f_ASAP7_75t_R EX___U767 ( .A(EX__n476), .Y(EX__n1572) );
  BUFx4f_ASAP7_75t_R EX___U768 ( .A(EX__n176), .Y(EX__n478) );
  BUFx6f_ASAP7_75t_R EX___U769 ( .A(forwarding_MEM_WB[25]), .Y(EX__n1492) );
  BUFx2_ASAP7_75t_R EX___U770 ( .A(EX__n864), .Y(EX__n479) );
  BUFx12f_ASAP7_75t_R EX___U771 ( .A(EX__n1258), .Y(EX__n480) );
  BUFx12f_ASAP7_75t_R EX___U772 ( .A(EX__n344), .Y(EX__n481) );
  BUFx12f_ASAP7_75t_R EX___U773 ( .A(EX__n1294), .Y(EX__n482) );
  BUFx4f_ASAP7_75t_R EX___U774 ( .A(EX__n484), .Y(EX__n483) );
  BUFx3_ASAP7_75t_R EX___U775 ( .A(EX__n438), .Y(EX__n484) );
  INVx4_ASAP7_75t_R EX___U776 ( .A(EX__n486), .Y(EX__n485) );
  BUFx12f_ASAP7_75t_R EX___U777 ( .A(EX__n487), .Y(EX__n486) );
  BUFx12f_ASAP7_75t_R EX___U778 ( .A(EX__n1572), .Y(EX__n487) );
  BUFx3_ASAP7_75t_R EX___U779 ( .A(EX__n489), .Y(EX__n488) );
  BUFx2_ASAP7_75t_R EX___U780 ( .A(input_data_2[22]), .Y(EX__n489) );
  BUFx16f_ASAP7_75t_R EX___U781 ( .A(EX__n736), .Y(EX__n490) );
  BUFx12f_ASAP7_75t_R EX___U782 ( .A(EX__n737), .Y(EX__n736) );
  BUFx2_ASAP7_75t_R EX___U783 ( .A(EX__n1433), .Y(EX__n491) );
  BUFx2_ASAP7_75t_R EX___U784 ( .A(EX__n1432), .Y(EX__n492) );
  CKINVDCx20_ASAP7_75t_R EX___U785 ( .A(EX__n1151), .Y(EX__n493) );
  CKINVDCx20_ASAP7_75t_R EX___U786 ( .A(EX__n493), .Y(EX__n494) );
  BUFx12f_ASAP7_75t_R EX___U787 ( .A(input_A[26]), .Y(EX__n495) );
  BUFx4f_ASAP7_75t_R EX___U788 ( .A(EX__n497), .Y(EX__n496) );
  BUFx3_ASAP7_75t_R EX___U789 ( .A(EX__n345), .Y(EX__n497) );
  BUFx4f_ASAP7_75t_R EX___U790 ( .A(EX__n499), .Y(EX__n498) );
  BUFx3_ASAP7_75t_R EX___U791 ( .A(EX__n346), .Y(EX__n499) );
  CKINVDCx20_ASAP7_75t_R EX___U792 ( .A(EX__n315), .Y(EX__n500) );
  CKINVDCx20_ASAP7_75t_R EX___U793 ( .A(EX__n500), .Y(EX__n501) );
  BUFx12_ASAP7_75t_R EX___U794 ( .A(input_data_2[3]), .Y(EX__n1186) );
  BUFx12f_ASAP7_75t_R EX___U795 ( .A(input_A[31]), .Y(EX__n503) );
  BUFx4f_ASAP7_75t_R EX___U796 ( .A(EX__n505), .Y(EX__n504) );
  BUFx3_ASAP7_75t_R EX___U797 ( .A(EX__n418), .Y(EX__n505) );
  BUFx4f_ASAP7_75t_R EX___U798 ( .A(EX__n507), .Y(EX__n506) );
  BUFx3_ASAP7_75t_R EX___U799 ( .A(EX__n419), .Y(EX__n507) );
  BUFx4f_ASAP7_75t_R EX___U800 ( .A(EX__n167), .Y(EX__n509) );
  BUFx2_ASAP7_75t_R EX___U801 ( .A(EX__n1042), .Y(EX__n510) );
  BUFx2_ASAP7_75t_R EX___U802 ( .A(EX__n670), .Y(EX__n511) );
  BUFx3_ASAP7_75t_R EX___U803 ( .A(EX__n559), .Y(EX__n915) );
  BUFx12f_ASAP7_75t_R EX___U804 ( .A(EX__n1354), .Y(EX__n514) );
  INVx2_ASAP7_75t_R EX___U805 ( .A(EX__n756), .Y(EX__n1336) );
  BUFx12f_ASAP7_75t_R EX___U806 ( .A(EX__n253), .Y(EX__n1340) );
  BUFx3_ASAP7_75t_R EX___U807 ( .A(EX__n516), .Y(EX__n515) );
  BUFx2_ASAP7_75t_R EX___U808 ( .A(EX__n1495), .Y(EX__n516) );
  BUFx12f_ASAP7_75t_R EX___U809 ( .A(EX__n519), .Y(EX__n517) );
  BUFx12f_ASAP7_75t_R EX___U810 ( .A(EX__n520), .Y(EX__n518) );
  BUFx12f_ASAP7_75t_R EX___U811 ( .A(EX__n267), .Y(EX__n519) );
  BUFx12f_ASAP7_75t_R EX___U812 ( .A(EX__n266), .Y(EX__n520) );
  BUFx12f_ASAP7_75t_R EX___U813 ( .A(EX__n759), .Y(EX__n1368) );
  BUFx3_ASAP7_75t_R EX___U814 ( .A(EX__n523), .Y(EX__n522) );
  BUFx2_ASAP7_75t_R EX___U815 ( .A(input_data_2[19]), .Y(EX__n523) );
  BUFx12f_ASAP7_75t_R EX___U816 ( .A(EX__n775), .Y(EX__n524) );
  BUFx4f_ASAP7_75t_R EX___U817 ( .A(EX__n522), .Y(EX__n776) );
  CKINVDCx20_ASAP7_75t_R EX___U818 ( .A(EX__n442), .Y(EX__n767) );
  CKINVDCx20_ASAP7_75t_R EX___U819 ( .A(EX__n1121), .Y(EX__n525) );
  BUFx16f_ASAP7_75t_R EX___U820 ( .A(EX__n1122), .Y(EX__n1121) );
  BUFx16f_ASAP7_75t_R EX___U821 ( .A(EX__n893), .Y(EX__n616) );
  INVx6_ASAP7_75t_R EX___U822 ( .A(EX__n660), .Y(EX__n893) );
  BUFx4f_ASAP7_75t_R EX___U823 ( .A(EX__n218), .Y(EX__n527) );
  BUFx3_ASAP7_75t_R EX___U824 ( .A(EX_read_reg_data_2[9]), .Y(EX__n1545) );
  BUFx2_ASAP7_75t_R EX___U825 ( .A(EX__n622), .Y(EX__n528) );
  BUFx2_ASAP7_75t_R EX___U826 ( .A(EX__n638), .Y(EX__n529) );
  BUFx3_ASAP7_75t_R EX___U827 ( .A(EX__n640), .Y(EX__n1047) );
  BUFx3_ASAP7_75t_R EX___U828 ( .A(EX__n535), .Y(EX__n534) );
  BUFx2_ASAP7_75t_R EX___U829 ( .A(EX__n1546), .Y(EX__n535) );
  BUFx3_ASAP7_75t_R EX___U830 ( .A(EX__n537), .Y(EX__n536) );
  BUFx2_ASAP7_75t_R EX___U831 ( .A(input_data_2[13]), .Y(EX__n537) );
  BUFx12f_ASAP7_75t_R EX___U832 ( .A(EX__n765), .Y(EX__n538) );
  BUFx4f_ASAP7_75t_R EX___U833 ( .A(EX__n536), .Y(EX__n766) );
  BUFx12f_ASAP7_75t_R EX___U834 ( .A(input_A[9]), .Y(EX__n539) );
  BUFx4f_ASAP7_75t_R EX___U835 ( .A(EX__n541), .Y(EX__n540) );
  BUFx3_ASAP7_75t_R EX___U836 ( .A(EX__n152), .Y(EX__n541) );
  BUFx4f_ASAP7_75t_R EX___U837 ( .A(EX__n543), .Y(EX__n542) );
  BUFx3_ASAP7_75t_R EX___U838 ( .A(EX__n153), .Y(EX__n543) );
  CKINVDCx20_ASAP7_75t_R EX___U839 ( .A(EX__n545), .Y(EX__n544) );
  BUFx16f_ASAP7_75t_R EX___U840 ( .A(EX__n1179), .Y(EX__n545) );
  BUFx12f_ASAP7_75t_R EX___U841 ( .A(EX__n894), .Y(EX__n660) );
  CKINVDCx16_ASAP7_75t_R EX___U842 ( .A(EX__n1251), .Y(EX__n778) );
  INVx13_ASAP7_75t_R EX___U843 ( .A(EX__n778), .Y(EX__n779) );
  CKINVDCx16_ASAP7_75t_R EX___U844 ( .A(EX__n470), .Y(EX__n547) );
  BUFx2_ASAP7_75t_R EX___U845 ( .A(input_data_2[16]), .Y(EX__n549) );
  BUFx4f_ASAP7_75t_R EX___U846 ( .A(EX__n204), .Y(EX__n551) );
  CKINVDCx11_ASAP7_75t_R EX___U847 ( .A(EX__n188), .Y(EX__n1164) );
  BUFx2_ASAP7_75t_R EX___U848 ( .A(EX__n994), .Y(EX__n554) );
  BUFx4f_ASAP7_75t_R EX___U849 ( .A(EX__n1492), .Y(EX__n555) );
  BUFx2_ASAP7_75t_R EX___U850 ( .A(EX__n1630), .Y(EX__n556) );
  INVx1_ASAP7_75t_R EX___U851 ( .A(EX__n915), .Y(EX__n558) );
  BUFx2_ASAP7_75t_R EX___U852 ( .A(EX__n560), .Y(EX__n559) );
  BUFx2_ASAP7_75t_R EX___U853 ( .A(EX__n1522), .Y(EX__n560) );
  BUFx3_ASAP7_75t_R EX___U854 ( .A(EX__n562), .Y(EX__n561) );
  BUFx2_ASAP7_75t_R EX___U855 ( .A(input_data_2[21]), .Y(EX__n562) );
  BUFx16f_ASAP7_75t_R EX___U856 ( .A(EX__n813), .Y(EX__n563) );
  BUFx12f_ASAP7_75t_R EX___U857 ( .A(EX__n814), .Y(EX__n813) );
  BUFx3_ASAP7_75t_R EX___U858 ( .A(EX__n565), .Y(EX__n564) );
  BUFx2_ASAP7_75t_R EX___U859 ( .A(input_data_2[5]), .Y(EX__n565) );
  BUFx16f_ASAP7_75t_R EX___U860 ( .A(EX__n1130), .Y(EX__n566) );
  BUFx12f_ASAP7_75t_R EX___U861 ( .A(EX__n797), .Y(EX__n796) );
  BUFx12f_ASAP7_75t_R EX___U862 ( .A(EX__n796), .Y(EX__n1130) );
  BUFx3_ASAP7_75t_R EX___U863 ( .A(EX__n568), .Y(EX__n567) );
  BUFx2_ASAP7_75t_R EX___U864 ( .A(EX__n1477), .Y(EX__n568) );
  BUFx3_ASAP7_75t_R EX___U865 ( .A(EX__n571), .Y(EX__n570) );
  BUFx2_ASAP7_75t_R EX___U866 ( .A(EX__n1498), .Y(EX__n571) );
  BUFx3_ASAP7_75t_R EX___U867 ( .A(EX__n413), .Y(EX__n573) );
  BUFx3_ASAP7_75t_R EX___U868 ( .A(EX__n575), .Y(EX__n574) );
  BUFx2_ASAP7_75t_R EX___U869 ( .A(EX__n1539), .Y(EX__n575) );
  BUFx3_ASAP7_75t_R EX___U870 ( .A(EX__n579), .Y(EX__n578) );
  BUFx2_ASAP7_75t_R EX___U871 ( .A(EX__n1564), .Y(EX__n579) );
  BUFx3_ASAP7_75t_R EX___U872 ( .A(EX__n583), .Y(EX__n582) );
  BUFx2_ASAP7_75t_R EX___U873 ( .A(EX__n1573), .Y(EX__n583) );
  BUFx2_ASAP7_75t_R EX___U874 ( .A(EX__n1445), .Y(EX__n585) );
  BUFx2_ASAP7_75t_R EX___U875 ( .A(EX__n1444), .Y(EX__n586) );
  CKINVDCx20_ASAP7_75t_R EX___U876 ( .A(EX__n1113), .Y(EX__n587) );
  CKINVDCx20_ASAP7_75t_R EX___U877 ( .A(EX__n587), .Y(EX__n588) );
  BUFx2_ASAP7_75t_R EX___U878 ( .A(input_data_2[25]), .Y(EX__n589) );
  BUFx12f_ASAP7_75t_R EX___U879 ( .A(EX__n591), .Y(EX__n590) );
  BUFx12f_ASAP7_75t_R EX___U880 ( .A(EX__n1157), .Y(EX__n591) );
  CKINVDCx14_ASAP7_75t_R EX___U881 ( .A(EX__n1156), .Y(EX__n592) );
  INVx6_ASAP7_75t_R EX___U882 ( .A(EX__n590), .Y(EX__n848) );
  BUFx16f_ASAP7_75t_R EX___U883 ( .A(EX__n848), .Y(EX__n1156) );
  BUFx12f_ASAP7_75t_R EX___U884 ( .A(EX__n661), .Y(EX__n1179) );
  BUFx12f_ASAP7_75t_R EX___U885 ( .A(input_A[30]), .Y(EX__n593) );
  BUFx4f_ASAP7_75t_R EX___U886 ( .A(EX__n595), .Y(EX__n594) );
  BUFx3_ASAP7_75t_R EX___U887 ( .A(EX__n392), .Y(EX__n595) );
  BUFx4f_ASAP7_75t_R EX___U888 ( .A(EX__n597), .Y(EX__n596) );
  BUFx3_ASAP7_75t_R EX___U889 ( .A(EX__n393), .Y(EX__n597) );
  BUFx12f_ASAP7_75t_R EX___U890 ( .A(input_A[4]), .Y(EX__n598) );
  CKINVDCx20_ASAP7_75t_R EX___U891 ( .A(EX__n1173), .Y(EX__n599) );
  CKINVDCx20_ASAP7_75t_R EX___U892 ( .A(EX__n599), .Y(EX__n600) );
  BUFx2_ASAP7_75t_R EX___U893 ( .A(EX__n1454), .Y(EX__n601) );
  BUFx2_ASAP7_75t_R EX___U894 ( .A(EX__n1453), .Y(EX__n602) );
  BUFx2_ASAP7_75t_R EX___U895 ( .A(EX__n1044), .Y(EX__n603) );
  BUFx2_ASAP7_75t_R EX___U896 ( .A(EX__n753), .Y(EX__n604) );
  BUFx12f_ASAP7_75t_R EX___U897 ( .A(EX__n324), .Y(EX__n605) );
  BUFx12f_ASAP7_75t_R EX___U898 ( .A(EX__n608), .Y(EX__n606) );
  BUFx12f_ASAP7_75t_R EX___U899 ( .A(EX__n1278), .Y(EX__n607) );
  BUFx12f_ASAP7_75t_R EX___U900 ( .A(EX__n323), .Y(EX__n608) );
  BUFx12f_ASAP7_75t_R EX___U901 ( .A(EX__n629), .Y(EX__n1278) );
  BUFx16f_ASAP7_75t_R EX___U902 ( .A(EX__n1106), .Y(EX__n609) );
  BUFx2_ASAP7_75t_R EX___U903 ( .A(EX__n1409), .Y(EX__n610) );
  BUFx2_ASAP7_75t_R EX___U904 ( .A(EX__n1408), .Y(EX__n611) );
  BUFx12f_ASAP7_75t_R EX___U905 ( .A(EX__n744), .Y(EX__n1106) );
  BUFx3_ASAP7_75t_R EX___U906 ( .A(EX__n613), .Y(EX__n612) );
  BUFx2_ASAP7_75t_R EX___U907 ( .A(input_data_2[20]), .Y(EX__n613) );
  BUFx12f_ASAP7_75t_R EX___U908 ( .A(EX__n699), .Y(EX__n614) );
  INVx6_ASAP7_75t_R EX___U909 ( .A(EX__n654), .Y(EX__n696) );
  BUFx16f_ASAP7_75t_R EX___U910 ( .A(EX__n1239), .Y(EX__n615) );
  CKINVDCx16_ASAP7_75t_R EX___U911 ( .A(EX__n615), .Y(EX__n1237) );
  BUFx12f_ASAP7_75t_R EX___U912 ( .A(EX__n634), .Y(EX__n1239) );
  BUFx10_ASAP7_75t_R EX___U913 ( .A(EX__n618), .Y(EX__n617) );
  BUFx4f_ASAP7_75t_R EX___U914 ( .A(EX__n228), .Y(EX__n618) );
  BUFx16f_ASAP7_75t_R EX___U915 ( .A(EX__n230), .Y(EX__n1077) );
  BUFx2_ASAP7_75t_R EX___U916 ( .A(EX__n1079), .Y(EX__n620) );
  BUFx2_ASAP7_75t_R EX___U917 ( .A(EX__n946), .Y(EX__n621) );
  CKINVDCx20_ASAP7_75t_R EX___U918 ( .A(EX__n1104), .Y(EX__n1105) );
  CKINVDCx14_ASAP7_75t_R EX___U919 ( .A(EX__n655), .Y(EX__n623) );
  BUFx12f_ASAP7_75t_R EX___U920 ( .A(EX__n697), .Y(EX__n654) );
  BUFx12f_ASAP7_75t_R EX___U921 ( .A(EX__n626), .Y(EX__n624) );
  BUFx12f_ASAP7_75t_R EX___U922 ( .A(EX__n342), .Y(EX__n625) );
  BUFx12f_ASAP7_75t_R EX___U923 ( .A(EX__n455), .Y(EX__n626) );
  BUFx12f_ASAP7_75t_R EX___U924 ( .A(EX__n1292), .Y(EX__n627) );
  BUFx12f_ASAP7_75t_R EX___U925 ( .A(EX__n1085), .Y(EX__n1292) );
  BUFx12f_ASAP7_75t_R EX___U926 ( .A(EX__n307), .Y(EX__n628) );
  BUFx12f_ASAP7_75t_R EX___U927 ( .A(EX__n306), .Y(EX__n629) );
  BUFx12f_ASAP7_75t_R EX___U928 ( .A(EX__n1275), .Y(EX__n1279) );
  BUFx12f_ASAP7_75t_R EX___U929 ( .A(EX__n631), .Y(EX__n630) );
  BUFx12f_ASAP7_75t_R EX___U930 ( .A(EX__n1261), .Y(EX__n631) );
  BUFx12f_ASAP7_75t_R EX___U931 ( .A(EX__n273), .Y(EX__n1261) );
  BUFx16f_ASAP7_75t_R EX___U932 ( .A(EX__n1244), .Y(EX__n632) );
  CKINVDCx16_ASAP7_75t_R EX___U933 ( .A(EX__n632), .Y(EX__n1242) );
  BUFx12f_ASAP7_75t_R EX___U934 ( .A(EX__n666), .Y(EX__n1244) );
  BUFx12f_ASAP7_75t_R EX___U935 ( .A(n50), .Y(EX__n633) );
  BUFx12f_ASAP7_75t_R EX___U936 ( .A(input_A[25]), .Y(EX__n634) );
  BUFx2_ASAP7_75t_R EX___U937 ( .A(EX__n1391), .Y(EX__n635) );
  BUFx2_ASAP7_75t_R EX___U938 ( .A(EX__n1390), .Y(EX__n636) );
  BUFx16f_ASAP7_75t_R EX___U939 ( .A(EX__n1250), .Y(EX__n1249) );
  INVx1_ASAP7_75t_R EX___U940 ( .A(EX__n735), .Y(EX__n638) );
  BUFx2_ASAP7_75t_R EX___U941 ( .A(EX__n641), .Y(EX__n640) );
  BUFx2_ASAP7_75t_R EX___U942 ( .A(EX__n1491), .Y(EX__n641) );
  CKINVDCx16_ASAP7_75t_R EX___U943 ( .A(EX__n687), .Y(EX__n1095) );
  BUFx3_ASAP7_75t_R EX___U944 ( .A(EX__n643), .Y(EX__n642) );
  BUFx2_ASAP7_75t_R EX___U945 ( .A(EX__n1524), .Y(EX__n643) );
  BUFx4f_ASAP7_75t_R EX___U946 ( .A(EX__n645), .Y(EX__n644) );
  BUFx3_ASAP7_75t_R EX___U947 ( .A(EX__n556), .Y(EX__n645) );
  BUFx3_ASAP7_75t_R EX___U948 ( .A(EX__n647), .Y(EX__n646) );
  BUFx2_ASAP7_75t_R EX___U949 ( .A(EX__n1531), .Y(EX__n647) );
  BUFx3_ASAP7_75t_R EX___U950 ( .A(EX__n649), .Y(EX__n648) );
  BUFx2_ASAP7_75t_R EX___U951 ( .A(input_data_2[24]), .Y(EX__n649) );
  BUFx12f_ASAP7_75t_R EX___U952 ( .A(EX__n953), .Y(EX__n650) );
  BUFx3_ASAP7_75t_R EX___U953 ( .A(EX__n652), .Y(EX__n651) );
  BUFx2_ASAP7_75t_R EX___U954 ( .A(input_data_2[14]), .Y(EX__n652) );
  BUFx12f_ASAP7_75t_R EX___U955 ( .A(EX__n792), .Y(EX__n653) );
  BUFx16f_ASAP7_75t_R EX___U956 ( .A(EX__n696), .Y(EX__n655) );
  BUFx12f_ASAP7_75t_R EX___U957 ( .A(EX__n698), .Y(EX__n697) );
  BUFx3_ASAP7_75t_R EX___U958 ( .A(EX__n658), .Y(EX__n657) );
  BUFx2_ASAP7_75t_R EX___U959 ( .A(EX__n1550), .Y(EX__n658) );
  BUFx3_ASAP7_75t_R EX___U960 ( .A(EX_read_reg_data_2[7]), .Y(EX__n659) );
  BUFx12f_ASAP7_75t_R EX___U961 ( .A(input_A[23]), .Y(EX__n661) );
  CKINVDCx20_ASAP7_75t_R EX___U962 ( .A(EX__n544), .Y(EX__n662) );
  CKINVDCx20_ASAP7_75t_R EX___U963 ( .A(EX__n662), .Y(EX__n663) );
  BUFx2_ASAP7_75t_R EX___U964 ( .A(EX__n1397), .Y(EX__n664) );
  BUFx2_ASAP7_75t_R EX___U965 ( .A(EX__n1396), .Y(EX__n665) );
  BUFx12f_ASAP7_75t_R EX___U966 ( .A(input_A[17]), .Y(EX__n666) );
  BUFx2_ASAP7_75t_R EX___U967 ( .A(EX__n1415), .Y(EX__n667) );
  BUFx2_ASAP7_75t_R EX___U968 ( .A(EX__n1414), .Y(EX__n668) );
  CKINVDCx16_ASAP7_75t_R EX___U969 ( .A(EX__n1242), .Y(EX__n1243) );
  INVx1_ASAP7_75t_R EX___U970 ( .A(EX__n1471), .Y(EX__n669) );
  BUFx3_ASAP7_75t_R EX___U971 ( .A(EX__n675), .Y(EX__n674) );
  BUFx2_ASAP7_75t_R EX___U972 ( .A(EX__n1563), .Y(EX__n675) );
  BUFx3_ASAP7_75t_R EX___U973 ( .A(EX__n678), .Y(EX__n677) );
  BUFx2_ASAP7_75t_R EX___U974 ( .A(EX__n1480), .Y(EX__n678) );
  BUFx3_ASAP7_75t_R EX___U975 ( .A(EX__n682), .Y(EX__n681) );
  BUFx2_ASAP7_75t_R EX___U976 ( .A(EX__n1501), .Y(EX__n682) );
  BUFx4f_ASAP7_75t_R EX___U977 ( .A(EX__n684), .Y(EX__n683) );
  BUFx3_ASAP7_75t_R EX___U978 ( .A(EX__n390), .Y(EX__n684) );
  BUFx3_ASAP7_75t_R EX___U979 ( .A(EX__n686), .Y(EX__n685) );
  BUFx2_ASAP7_75t_R EX___U980 ( .A(EX__n1543), .Y(EX__n686) );
  BUFx16f_ASAP7_75t_R EX___U981 ( .A(EX__n1097), .Y(EX__n687) );
  BUFx2_ASAP7_75t_R EX___U982 ( .A(EX__n1459), .Y(EX__n688) );
  BUFx2_ASAP7_75t_R EX___U983 ( .A(EX__n1460), .Y(EX__n689) );
  BUFx12f_ASAP7_75t_R EX___U984 ( .A(EX__n739), .Y(EX__n1097) );
  BUFx4f_ASAP7_75t_R EX___U985 ( .A(EX__n691), .Y(EX__n690) );
  BUFx3_ASAP7_75t_R EX___U986 ( .A(EX__n6), .Y(EX__EX__n691) );
  BUFx3_ASAP7_75t_R EX___U987 ( .A(EX__n693), .Y(EX__n692) );
  BUFx2_ASAP7_75t_R EX___U988 ( .A(EX__n1568), .Y(EX__n693) );
  INVx1_ASAP7_75t_R EX___U989 ( .A(EX__n1203), .Y(EX_read_reg_data_2[1]) );
  BUFx12f_ASAP7_75t_R EX___U990 ( .A(EX__n889), .Y(EX__n698) );
  BUFx10_ASAP7_75t_R EX___U991 ( .A(input_data_2[31]), .Y(EX__n889) );
  BUFx10_ASAP7_75t_R EX___U992 ( .A(EX__n700), .Y(EX__n699) );
  BUFx4f_ASAP7_75t_R EX___U993 ( .A(EX__n612), .Y(EX__n700) );
  BUFx16f_ASAP7_75t_R EX___U994 ( .A(EX__n614), .Y(EX__n1031) );
  BUFx2_ASAP7_75t_R EX___U995 ( .A(EX__n1082), .Y(EX__n702) );
  BUFx2_ASAP7_75t_R EX___U996 ( .A(EX__n996), .Y(EX__n703) );
  BUFx3_ASAP7_75t_R EX___U997 ( .A(EX__n876), .Y(EX__n875) );
  BUFx3_ASAP7_75t_R EX___U998 ( .A(EX__n708), .Y(EX__n707) );
  BUFx2_ASAP7_75t_R EX___U999 ( .A(EX__n1470), .Y(EX__n708) );
  BUFx3_ASAP7_75t_R EX___U1000 ( .A(EX__n712), .Y(EX__n711) );
  BUFx2_ASAP7_75t_R EX___U1001 ( .A(EX__n1515), .Y(EX__n712) );
  BUFx3_ASAP7_75t_R EX___U1002 ( .A(EX__n714), .Y(EX__n713) );
  BUFx2_ASAP7_75t_R EX___U1003 ( .A(input_data_2[23]), .Y(EX__n714) );
  BUFx12f_ASAP7_75t_R EX___U1004 ( .A(EX__n1054), .Y(EX__n715) );
  BUFx3_ASAP7_75t_R EX___U1005 ( .A(EX__n411), .Y(EX__n717) );
  BUFx3_ASAP7_75t_R EX___U1006 ( .A(EX__n719), .Y(EX__n718) );
  BUFx2_ASAP7_75t_R EX___U1007 ( .A(EX__n1484), .Y(EX__n719) );
  BUFx3_ASAP7_75t_R EX___U1008 ( .A(EX_read_reg_data_2[27]), .Y(EX__n720) );
  INVx2_ASAP7_75t_R EX___U1009 ( .A(EX__n716), .Y(EX_read_reg_data_2[27]) );
  BUFx3_ASAP7_75t_R EX___U1010 ( .A(EX__n724), .Y(EX__n723) );
  BUFx2_ASAP7_75t_R EX___U1011 ( .A(EX__n1536), .Y(EX__n724) );
  BUFx3_ASAP7_75t_R EX___U1012 ( .A(EX__n728), .Y(EX__n727) );
  BUFx2_ASAP7_75t_R EX___U1013 ( .A(EX__n1554), .Y(EX__n728) );
  BUFx3_ASAP7_75t_R EX___U1014 ( .A(EX__n730), .Y(EX__n1541) );
  INVx1_ASAP7_75t_R EX___U1015 ( .A(EX__n555), .Y(EX__n734) );
  BUFx4f_ASAP7_75t_R EX___U1016 ( .A(EX__n488), .Y(EX__n737) );
  BUFx2_ASAP7_75t_R EX___U1017 ( .A(EX__n1163), .Y(EX__n738) );
  BUFx12f_ASAP7_75t_R EX___U1018 ( .A(input_A[2]), .Y(EX__n739) );
  BUFx4f_ASAP7_75t_R EX___U1019 ( .A(EX__n741), .Y(EX__n740) );
  BUFx3_ASAP7_75t_R EX___U1020 ( .A(EX__n689), .Y(EX__n741) );
  BUFx4f_ASAP7_75t_R EX___U1021 ( .A(EX__n743), .Y(EX__n742) );
  BUFx3_ASAP7_75t_R EX___U1022 ( .A(EX__n688), .Y(EX__n743) );
  INVx2_ASAP7_75t_R EX___U1023 ( .A(EX__n1340), .Y(EX__n1335) );
  CKINVDCx16_ASAP7_75t_R EX___U1024 ( .A(EX__n1095), .Y(EX__n1096) );
  BUFx12f_ASAP7_75t_R EX___U1025 ( .A(input_A[19]), .Y(EX__n744) );
  BUFx4f_ASAP7_75t_R EX___U1026 ( .A(EX__n746), .Y(EX__n745) );
  BUFx3_ASAP7_75t_R EX___U1027 ( .A(EX__n610), .Y(EX__n746) );
  BUFx4f_ASAP7_75t_R EX___U1028 ( .A(EX__n748), .Y(EX__n747) );
  BUFx3_ASAP7_75t_R EX___U1029 ( .A(EX__n611), .Y(EX__n748) );
  CKINVDCx20_ASAP7_75t_R EX___U1030 ( .A(EX__n525), .Y(EX__n749) );
  BUFx12f_ASAP7_75t_R EX___U1031 ( .A(EX__n751), .Y(EX__n750) );
  BUFx12f_ASAP7_75t_R EX___U1032 ( .A(input_data_2[1]), .Y(EX__n751) );
  INVx6_ASAP7_75t_R EX___U1033 ( .A(EX__n750), .Y(EX__n1122) );
  BUFx2_ASAP7_75t_R EX___U1034 ( .A(EX__n995), .Y(EX__n752) );
  INVx1_ASAP7_75t_R EX___U1035 ( .A(EX__n908), .Y(EX__n753) );
  BUFx12f_ASAP7_75t_R EX___U1036 ( .A(EX__n756), .Y(EX__n754) );
  BUFx12f_ASAP7_75t_R EX___U1037 ( .A(EX__n269), .Y(EX__n756) );
  BUFx12f_ASAP7_75t_R EX___U1038 ( .A(EX__n268), .Y(EX__n757) );
  BUFx12f_ASAP7_75t_R EX___U1039 ( .A(EX__n1337), .Y(EX__n1338) );
  BUFx10_ASAP7_75t_R EX___U1040 ( .A(EX__n139), .Y(EX__n1355) );
  BUFx12f_ASAP7_75t_R EX___U1041 ( .A(EX__n401), .Y(EX__n758) );
  BUFx12f_ASAP7_75t_R EX___U1042 ( .A(EX__n401), .Y(EX__n759) );
  BUFx12f_ASAP7_75t_R EX___U1043 ( .A(EX__n1365), .Y(EX__n1369) );
  BUFx12f_ASAP7_75t_R EX___U1044 ( .A(EX__n1291), .Y(EX__n760) );
  BUFx12f_ASAP7_75t_R EX___U1045 ( .A(EX__n624), .Y(EX__n1291) );
  INVx2_ASAP7_75t_R EX___U1046 ( .A(ID_EX_imm[19]), .Y(EX__n1514) );
  BUFx6f_ASAP7_75t_R EX___U1047 ( .A(EX__n1280), .Y(EX__n1269) );
  BUFx6f_ASAP7_75t_R EX___U1048 ( .A(EX__n1266), .Y(EX__n1268) );
  BUFx6f_ASAP7_75t_R EX___U1049 ( .A(EX__n1265), .Y(EX__n1267) );
  BUFx12f_ASAP7_75t_R EX___U1050 ( .A(EX__n1260), .Y(EX__n761) );
  BUFx12f_ASAP7_75t_R EX___U1051 ( .A(EX__n1262), .Y(EX__n1260) );
  BUFx2_ASAP7_75t_R EX___U1052 ( .A(EX__n1117), .Y(EX__n764) );
  BUFx6f_ASAP7_75t_R EX___U1053 ( .A(EX__n766), .Y(EX__n765) );
  INVx1_ASAP7_75t_R EX___U1054 ( .A(EX__n1533), .Y(EX__n1117) );
  BUFx2_ASAP7_75t_R EX___U1055 ( .A(EX__n804), .Y(EX__n768) );
  BUFx2_ASAP7_75t_R EX___U1056 ( .A(EX__n806), .Y(EX__n769) );
  BUFx12f_ASAP7_75t_R EX___U1057 ( .A(input_A[7]), .Y(EX__n770) );
  BUFx4f_ASAP7_75t_R EX___U1058 ( .A(EX__n772), .Y(EX__n771) );
  BUFx3_ASAP7_75t_R EX___U1059 ( .A(EX__n585), .Y(EX__n772) );
  BUFx4f_ASAP7_75t_R EX___U1060 ( .A(EX__n774), .Y(EX__n773) );
  BUFx3_ASAP7_75t_R EX___U1061 ( .A(EX__n586), .Y(EX__n774) );
  BUFx6f_ASAP7_75t_R EX___U1062 ( .A(EX__n1289), .Y(EX__n1287) );
  BUFx12f_ASAP7_75t_R EX___U1063 ( .A(EX__n1293), .Y(EX__n1289) );
  BUFx6f_ASAP7_75t_R EX___U1064 ( .A(EX__n1277), .Y(EX__n1272) );
  BUFx6f_ASAP7_75t_R EX___U1065 ( .A(EX__n1277), .Y(EX__n1271) );
  BUFx6f_ASAP7_75t_R EX___U1066 ( .A(EX__n1277), .Y(EX__n1270) );
  BUFx12f_ASAP7_75t_R EX___U1067 ( .A(EX__n628), .Y(EX__n1277) );
  BUFx12f_ASAP7_75t_R EX___U1068 ( .A(EX__n630), .Y(EX__n1259) );
  BUFx12f_ASAP7_75t_R EX___U1069 ( .A(EX__n1370), .Y(EX__n1366) );
  BUFx6f_ASAP7_75t_R EX___U1070 ( .A(EX__n776), .Y(EX__n775) );
  CKINVDCx14_ASAP7_75t_R EX___U1071 ( .A(EX__n563), .Y(EX__n1075) );
  BUFx4f_ASAP7_75t_R EX___U1072 ( .A(EX__n729), .Y(EX__n1557) );
  INVx2_ASAP7_75t_R EX___U1073 ( .A(EX__n1557), .Y(EX__n780) );
  OA22x2_ASAP7_75t_R EX___U1074 ( .A1(EX__n780), .A2(EX__n1320), .B1(EX__n1556), .B2(EX__n1302), 
        .Y(input_data_2[6]) );
  BUFx2_ASAP7_75t_R EX___U1075 ( .A(EX__n805), .Y(EX__n783) );
  BUFx2_ASAP7_75t_R EX___U1076 ( .A(EX__n998), .Y(EX__n784) );
  BUFx6f_ASAP7_75t_R EX___U1077 ( .A(EX__n1352), .Y(EX__n1347) );
  BUFx6f_ASAP7_75t_R EX___U1078 ( .A(EX__n1352), .Y(EX__n1346) );
  BUFx6f_ASAP7_75t_R EX___U1079 ( .A(EX__n1352), .Y(EX__n1345) );
  BUFx12f_ASAP7_75t_R EX___U1080 ( .A(EX__n263), .Y(EX__n1352) );
  INVx2_ASAP7_75t_R EX___U1081 ( .A(EX__n1338), .Y(EX__n1326) );
  INVx2_ASAP7_75t_R EX___U1082 ( .A(EX__n1337), .Y(EX__n1327) );
  INVx2_ASAP7_75t_R EX___U1083 ( .A(EX__n1342), .Y(EX__n1328) );
  BUFx6f_ASAP7_75t_R EX___U1084 ( .A(ID_EX_imm[18]), .Y(EX__n786) );
  BUFx2_ASAP7_75t_R EX___U1085 ( .A(ID_EX_imm[18]), .Y(EX__n787) );
  BUFx6f_ASAP7_75t_R EX___U1086 ( .A(EX__n343), .Y(EX__n1286) );
  BUFx6f_ASAP7_75t_R EX___U1087 ( .A(EX__n455), .Y(EX__n1285) );
  BUFx6f_ASAP7_75t_R EX___U1088 ( .A(EX__n1291), .Y(EX__n1284) );
  BUFx12f_ASAP7_75t_R EX___U1089 ( .A(EX__n1280), .Y(EX__n1276) );
  BUFx6f_ASAP7_75t_R EX___U1090 ( .A(EX__n606), .Y(EX__n1274) );
  BUFx6f_ASAP7_75t_R EX___U1091 ( .A(EX__n1276), .Y(EX__n1273) );
  BUFx12f_ASAP7_75t_R EX___U1092 ( .A(EX__n273), .Y(EX__n1258) );
  BUFx6f_ASAP7_75t_R EX___U1093 ( .A(EX__n1370), .Y(EX__n1360) );
  BUFx6f_ASAP7_75t_R EX___U1094 ( .A(EX__n1357), .Y(EX__n1359) );
  BUFx10_ASAP7_75t_R EX___U1095 ( .A(EX__n789), .Y(EX__n788) );
  BUFx4f_ASAP7_75t_R EX___U1096 ( .A(EX__n443), .Y(EX__n789) );
  BUFx16f_ASAP7_75t_R EX___U1097 ( .A(EX__n445), .Y(EX__n1127) );
  CKINVDCx20_ASAP7_75t_R EX___U1098 ( .A(EX__n1127), .Y(EX__n790) );
  BUFx2_ASAP7_75t_R EX___U1099 ( .A(EX__n1129), .Y(EX__n791) );
  BUFx10_ASAP7_75t_R EX___U1100 ( .A(EX__n793), .Y(EX__n792) );
  BUFx4f_ASAP7_75t_R EX___U1101 ( .A(EX__n651), .Y(EX__n793) );
  BUFx16f_ASAP7_75t_R EX___U1102 ( .A(EX__n653), .Y(EX__n1170) );
  BUFx2_ASAP7_75t_R EX___U1103 ( .A(EX__n1172), .Y(EX__n795) );
  BUFx4f_ASAP7_75t_R EX___U1104 ( .A(EX__n564), .Y(EX__n797) );
  BUFx2_ASAP7_75t_R EX___U1105 ( .A(EX__n1131), .Y(EX__n799) );
  BUFx6f_ASAP7_75t_R EX___U1106 ( .A(ID_EX_imm[11]), .Y(EX__n1537) );
  INVx3_ASAP7_75t_R EX___U1107 ( .A(EX__n1537), .Y(EX__n800) );
  BUFx4f_ASAP7_75t_R EX___U1108 ( .A(EX__n726), .Y(EX__n1538) );
  INVx2_ASAP7_75t_R EX___U1109 ( .A(EX__n1538), .Y(EX__n801) );
  OA22x2_ASAP7_75t_R EX___U1110 ( .A1(EX__n801), .A2(EX__n1313), .B1(EX__n1300), .B2(EX__n800), .Y(
        input_data_2[11]) );
  BUFx2_ASAP7_75t_R EX___U1111 ( .A(EX__n980), .Y(EX__n803) );
  INVx1_ASAP7_75t_R EX___U1112 ( .A(EX__n945), .Y(EX__n806) );
  BUFx2_ASAP7_75t_R EX___U1113 ( .A(EX__n1641), .Y(EX__n807) );
  BUFx12f_ASAP7_75t_R EX___U1114 ( .A(EX__n289), .Y(EX__n1351) );
  BUFx12f_ASAP7_75t_R EX___U1115 ( .A(EX__n1355), .Y(EX__n1354) );
  BUFx6f_ASAP7_75t_R EX___U1116 ( .A(EX__n1367), .Y(EX__n1363) );
  BUFx6f_ASAP7_75t_R EX___U1117 ( .A(EX__n1367), .Y(EX__n1362) );
  BUFx6f_ASAP7_75t_R EX___U1118 ( .A(EX__n1367), .Y(EX__n1361) );
  BUFx12f_ASAP7_75t_R EX___U1119 ( .A(EX__n758), .Y(EX__n1367) );
  BUFx12f_ASAP7_75t_R EX___U1120 ( .A(EX__n423), .Y(EX__n1264) );
  INVx2_ASAP7_75t_R EX___U1121 ( .A(EX__n1339), .Y(EX__n1323) );
  INVx2_ASAP7_75t_R EX___U1122 ( .A(EX__n1339), .Y(EX__n1322) );
  INVx2_ASAP7_75t_R EX___U1123 ( .A(EX__n1339), .Y(EX__n1324) );
  BUFx12f_ASAP7_75t_R EX___U1124 ( .A(EX__n1340), .Y(EX__n1339) );
  INVx3_ASAP7_75t_R EX___U1125 ( .A(EX__n755), .Y(EX__n1325) );
  BUFx4f_ASAP7_75t_R EX___U1126 ( .A(EX__n439), .Y(EX__n810) );
  BUFx2_ASAP7_75t_R EX___U1127 ( .A(EX__n1223), .Y(EX__n811) );
  BUFx2_ASAP7_75t_R EX___U1128 ( .A(EX__n1224), .Y(EX__n812) );
  BUFx4f_ASAP7_75t_R EX___U1129 ( .A(EX__n561), .Y(EX__n814) );
  BUFx12f_ASAP7_75t_R EX___U1130 ( .A(EX__n816), .Y(EX__n815) );
  BUFx12f_ASAP7_75t_R EX___U1131 ( .A(input_data_2[2]), .Y(EX__n816) );
  BUFx2_ASAP7_75t_R EX___U1132 ( .A(EX__n1253), .Y(EX__n817) );
  BUFx2_ASAP7_75t_R EX___U1133 ( .A(EX__n1254), .Y(EX__n818) );
  BUFx16f_ASAP7_75t_R EX___U1134 ( .A(EX__n1252), .Y(EX__n1251) );
  INVx6_ASAP7_75t_R EX___U1135 ( .A(EX__n815), .Y(EX__n1252) );
  BUFx6f_ASAP7_75t_R EX___U1136 ( .A(ID_EX_imm[7]), .Y(EX__n1552) );
  INVx3_ASAP7_75t_R EX___U1137 ( .A(EX__n1552), .Y(EX__n819) );
  BUFx4f_ASAP7_75t_R EX___U1138 ( .A(EX__n659), .Y(EX__n1553) );
  INVx2_ASAP7_75t_R EX___U1139 ( .A(EX__n1553), .Y(EX__n820) );
  OA22x2_ASAP7_75t_R EX___U1140 ( .A1(EX__n820), .A2(EX__n1316), .B1(EX__n819), .B2(EX__n1302), .Y(
        input_data_2[7]) );
  BUFx3_ASAP7_75t_R EX___U1141 ( .A(EX__n829), .Y(EX__n828) );
  BUFx2_ASAP7_75t_R EX___U1142 ( .A(EX__n1474), .Y(EX__n829) );
  BUFx4f_ASAP7_75t_R EX___U1143 ( .A(EX__n831), .Y(EX__n830) );
  BUFx3_ASAP7_75t_R EX___U1144 ( .A(EX__n833), .Y(EX__n832) );
  BUFx2_ASAP7_75t_R EX___U1145 ( .A(EX__n1487), .Y(EX__n833) );
  BUFx3_ASAP7_75t_R EX___U1146 ( .A(EX__n837), .Y(EX__n836) );
  BUFx2_ASAP7_75t_R EX___U1147 ( .A(EX__n1509), .Y(EX__n837) );
  BUFx3_ASAP7_75t_R EX___U1148 ( .A(EX__n841), .Y(EX__n840) );
  BUFx2_ASAP7_75t_R EX___U1149 ( .A(EX__n1528), .Y(EX__n841) );
  BUFx12f_ASAP7_75t_R EX___U1150 ( .A(input_A[11]), .Y(EX__n843) );
  BUFx4f_ASAP7_75t_R EX___U1151 ( .A(EX__n845), .Y(EX__n844) );
  BUFx3_ASAP7_75t_R EX___U1152 ( .A(EX__n491), .Y(EX__n845) );
  BUFx4f_ASAP7_75t_R EX___U1153 ( .A(EX__n847), .Y(EX__n846) );
  BUFx3_ASAP7_75t_R EX___U1154 ( .A(EX__n492), .Y(EX__n847) );
  BUFx6f_ASAP7_75t_R EX___U1155 ( .A(EX__n849), .Y(EX__n1157) );
  BUFx4f_ASAP7_75t_R EX___U1156 ( .A(EX__n850), .Y(EX__n849) );
  BUFx3_ASAP7_75t_R EX___U1157 ( .A(EX__n589), .Y(EX__n850) );
  CKINVDCx16_ASAP7_75t_R EX___U1158 ( .A(EX__n592), .Y(EX__n851) );
  BUFx4f_ASAP7_75t_R EX___U1159 ( .A(ID_EX_imm[25]), .Y(EX__n1493) );
  OA21x2_ASAP7_75t_R EX___U1160 ( .A1(EX__n1283), .A2(EX__n62), .B(EX__n853), .Y(EX__n1633) );
  AO22x2_ASAP7_75t_R EX___U1161 ( .A1(forwarding_EX_MEM[10]), .A2(EX__n1272), .B1(
        ID_EX_read_reg_data_2[10]), .B2(EX__n1256), .Y(EX__n1539) );
  INVx1_ASAP7_75t_R EX___U1162 ( .A(EX__n574), .Y(EX__n853) );
  AO22x2_ASAP7_75t_R EX___U1163 ( .A1(forwarding_EX_MEM[2]), .A2(EX__n1274), .B1(
        ID_EX_read_reg_data_2[2]), .B2(EX__n457), .Y(EX__n1564) );
  INVx1_ASAP7_75t_R EX___U1164 ( .A(EX__n578), .Y(EX__n855) );
  BUFx10_ASAP7_75t_R EX___U1165 ( .A(EX__n857), .Y(EX__n856) );
  BUFx4f_ASAP7_75t_R EX___U1166 ( .A(EX__n424), .Y(EX__n857) );
  BUFx16f_ASAP7_75t_R EX___U1167 ( .A(EX__n426), .Y(EX__n1219) );
  BUFx2_ASAP7_75t_R EX___U1168 ( .A(EX__n1221), .Y(EX__n859) );
  OA22x2_ASAP7_75t_R EX___U1169 ( .A1(EX__n860), .A2(EX__n1313), .B1(EX__n1300), .B2(EX__n1535), 
        .Y(input_data_2[12]) );
  INVx1_ASAP7_75t_R EX___U1170 ( .A(EX__n913), .Y(EX_read_reg_data_2[16]) );
  INVx1_ASAP7_75t_R EX___U1171 ( .A(EX__n1083), .Y(EX__n864) );
  BUFx2_ASAP7_75t_R EX___U1172 ( .A(EX__n1191), .Y(EX__n881) );
  BUFx12f_ASAP7_75t_R EX___U1173 ( .A(EX__n625), .Y(EX__n1290) );
  BUFx12f_ASAP7_75t_R EX___U1174 ( .A(EX__n255), .Y(EX__n1353) );
  BUFx3_ASAP7_75t_R EX___U1175 ( .A(EX__n787), .Y(EX__n1516) );
  BUFx12f_ASAP7_75t_R EX___U1176 ( .A(EX__n757), .Y(EX__n885) );
  BUFx12f_ASAP7_75t_R EX___U1177 ( .A(EX__n754), .Y(EX__n886) );
  INVx2_ASAP7_75t_R EX___U1178 ( .A(EX__n886), .Y(EX__n1331) );
  INVx2_ASAP7_75t_R EX___U1179 ( .A(EX__n886), .Y(EX__n1330) );
  INVx2_ASAP7_75t_R EX___U1180 ( .A(EX__n886), .Y(EX__n1329) );
  CKINVDCx8_ASAP7_75t_R EX___U1181 ( .A(EX__n81), .Y(EX__n1332) );
  AND2x2_ASAP7_75t_R EX___U1182 ( .A(ForwardB[1]), .B(EX__n1468), .Y(EX__n1469) );
  BUFx12f_ASAP7_75t_R EX___U1183 ( .A(EX__n462), .Y(EX__n1370) );
  CKINVDCx16_ASAP7_75t_R EX___U1184 ( .A(EX__n623), .Y(EX__n888) );
  BUFx2_ASAP7_75t_R EX___U1185 ( .A(EX__n1248), .Y(EX__n890) );
  BUFx3_ASAP7_75t_R EX___U1186 ( .A(ID_EX_imm[31]), .Y(EX__n1472) );
  CKINVDCx20_ASAP7_75t_R EX___U1187 ( .A(EX__n616), .Y(EX__n891) );
  CKINVDCx20_ASAP7_75t_R EX___U1188 ( .A(EX__n891), .Y(EX__n892) );
  BUFx12f_ASAP7_75t_R EX___U1189 ( .A(EX__n895), .Y(EX__n894) );
  BUFx12f_ASAP7_75t_R EX___U1190 ( .A(input_data_2[0]), .Y(EX__n895) );
  BUFx2_ASAP7_75t_R EX___U1191 ( .A(EX__n1188), .Y(EX__n896) );
  BUFx3_ASAP7_75t_R EX___U1192 ( .A(EX__n732), .Y(EX__n1576) );
  OA22x2_ASAP7_75t_R EX___U1193 ( .A1(EX__n897), .A2(EX__n1312), .B1(EX__n1298), .B2(EX__n1514), 
        .Y(input_data_2[19]) );
  INVx2_ASAP7_75t_R EX___U1194 ( .A(EX__n1485), .Y(EX__n899) );
  BUFx4f_ASAP7_75t_R EX___U1195 ( .A(EX__n720), .Y(EX__n1486) );
  INVx2_ASAP7_75t_R EX___U1196 ( .A(EX__n1486), .Y(EX__n900) );
  OA22x2_ASAP7_75t_R EX___U1197 ( .A1(EX__n900), .A2(EX__n395), .B1(EX__n1295), .B2(EX__n899), .Y(
        input_data_2[27]) );
  BUFx3_ASAP7_75t_R EX___U1198 ( .A(EX__n907), .Y(EX__n906) );
  BUFx2_ASAP7_75t_R EX___U1199 ( .A(EX__n1505), .Y(EX__n907) );
  BUFx12f_ASAP7_75t_R EX___U1200 ( .A(ID_EX_ALUSrc), .Y(EX__n1321) );
  OA21x2_ASAP7_75t_R EX___U1201 ( .A1(EX__n626), .A2(EX__n1133), .B(EX__n910), .Y(EX__n1619) );
  AO22x2_ASAP7_75t_R EX___U1202 ( .A1(forwarding_EX_MEM[24]), .A2(EX__n1267), .B1(
        ID_EX_read_reg_data_2[24]), .B2(EX__n1256), .Y(EX__n1495) );
  INVx1_ASAP7_75t_R EX___U1203 ( .A(EX__n515), .Y(EX__n910) );
  OA21x2_ASAP7_75t_R EX___U1204 ( .A1(EX__n1285), .A2(EX__n882), .B(EX__n912), .Y(EX__n1625) );
  AO22x2_ASAP7_75t_R EX___U1205 ( .A1(forwarding_EX_MEM[18]), .A2(EX__n1269), .B1(
        ID_EX_read_reg_data_2[18]), .B2(EX__n1255), .Y(EX__n1515) );
  INVx1_ASAP7_75t_R EX___U1206 ( .A(EX__n711), .Y(EX__n912) );
  OA21x2_ASAP7_75t_R EX___U1207 ( .A1(EX__n1284), .A2(EX__n733), .B(EX__n558), .Y(EX__n1627) );
  AO22x2_ASAP7_75t_R EX___U1208 ( .A1(forwarding_EX_MEM[16]), .A2(EX__n1270), .B1(
        ID_EX_read_reg_data_2[16]), .B2(EX__n314), .Y(EX__n1522) );
  AO22x2_ASAP7_75t_R EX___U1209 ( .A1(forwarding_EX_MEM[0]), .A2(EX__n1275), .B1(
        ID_EX_read_reg_data_2[0]), .B2(EX__n1257), .Y(EX__n1573) );
  INVx1_ASAP7_75t_R EX___U1210 ( .A(EX__n582), .Y(EX__n917) );
  AO22x2_ASAP7_75t_R EX___U1211 ( .A1(EX__n763), .A2(ID_EX_ALUSrc), .B1(
        EX_read_reg_data_2[3]), .B2(EX__n1579), .Y(input_data_2[3]) );
  OR2x2_ASAP7_75t_R EX___U1212 ( .A(EX__n1333), .B(EX__n1380), .Y(EX__n1382) );
  INVx2_ASAP7_75t_R EX___U1213 ( .A(EX__n247), .Y(EX__n918) );
  OA22x2_ASAP7_75t_R EX___U1214 ( .A1(EX__n884), .A2(EX__n1357), .B1(EX__n1583), .B2(EX__n1354), 
        .Y(EX__n1381) );
  INVx2_ASAP7_75t_R EX___U1215 ( .A(EX__n249), .Y(EX__n919) );
  CKINVDCx20_ASAP7_75t_R EX___U1216 ( .A(EX__n252), .Y(EX__n920) );
  OR2x2_ASAP7_75t_R EX___U1217 ( .A(EX__n1329), .B(EX__n1419), .Y(EX__n1421) );
  INVx2_ASAP7_75t_R EX___U1218 ( .A(EX__n144), .Y(EX__n922) );
  OA22x2_ASAP7_75t_R EX___U1219 ( .A1(EX__n1361), .A2(EX__n621), .B1(EX__n1596), .B2(EX__n1348), 
        .Y(EX__n1420) );
  INVx2_ASAP7_75t_R EX___U1220 ( .A(EX__n146), .Y(EX__n923) );
  CKINVDCx20_ASAP7_75t_R EX___U1221 ( .A(EX__n88), .Y(EX__n924) );
  CKINVDCx20_ASAP7_75t_R EX___U1222 ( .A(EX__n924), .Y(EX__n925) );
  OR2x2_ASAP7_75t_R EX___U1223 ( .A(EX__n1332), .B(EX__n1440), .Y(EX__n1442) );
  INVx2_ASAP7_75t_R EX___U1224 ( .A(EX__n198), .Y(EX__n927) );
  OA22x2_ASAP7_75t_R EX___U1225 ( .A1(EX__n1363), .A2(EX__n703), .B1(EX__n1603), .B2(EX__n256), .Y(
        n1441) );
  INVx2_ASAP7_75t_R EX___U1226 ( .A(EX__n200), .Y(EX__n928) );
  CKINVDCx20_ASAP7_75t_R EX___U1227 ( .A(EX__n203), .Y(EX__n929) );
  BUFx3_ASAP7_75t_R EX___U1228 ( .A(EX__n826), .Y(EX__n932) );
  BUFx3_ASAP7_75t_R EX___U1229 ( .A(EX__n934), .Y(EX__n933) );
  BUFx2_ASAP7_75t_R EX___U1230 ( .A(EX__n1518), .Y(EX__n934) );
  BUFx3_ASAP7_75t_R EX___U1231 ( .A(EX__n938), .Y(EX__n937) );
  BUFx2_ASAP7_75t_R EX___U1232 ( .A(EX__n1534), .Y(EX__n938) );
  BUFx3_ASAP7_75t_R EX___U1233 ( .A(EX__n942), .Y(EX__n941) );
  BUFx2_ASAP7_75t_R EX___U1234 ( .A(EX__n1558), .Y(EX__n942) );
  BUFx3_ASAP7_75t_R EX___U1235 ( .A(ID_EX_imm[17]), .Y(EX__n1520) );
  INVx1_ASAP7_75t_R EX___U1236 ( .A(EX__n877), .Y(EX__n946) );
  OA21x2_ASAP7_75t_R EX___U1237 ( .A1(EX__n1287), .A2(EX__n989), .B(EX__n948), .Y(EX__n1614) );
  AO22x2_ASAP7_75t_R EX___U1238 ( .A1(forwarding_EX_MEM[29]), .A2(EX__n1265), .B1(
        ID_EX_read_reg_data_2[29]), .B2(EX__n1261), .Y(EX__n1477) );
  INVx1_ASAP7_75t_R EX___U1239 ( .A(EX__n567), .Y(EX__n948) );
  AO22x2_ASAP7_75t_R EX___U1240 ( .A1(forwarding_EX_MEM[20]), .A2(EX__n1268), .B1(
        ID_EX_read_reg_data_2[20]), .B2(EX__n270), .Y(EX__n1509) );
  INVx1_ASAP7_75t_R EX___U1241 ( .A(EX__n836), .Y(EX__n950) );
  OA21x2_ASAP7_75t_R EX___U1242 ( .A1(EX__n1282), .A2(EX__n1040), .B(EX__n952), .Y(EX__n1634) );
  INVx2_ASAP7_75t_R EX___U1243 ( .A(EX__n683), .Y(EX_read_reg_data_2[9]) );
  AO22x2_ASAP7_75t_R EX___U1244 ( .A1(forwarding_EX_MEM[9]), .A2(EX__n1272), .B1(
        ID_EX_read_reg_data_2[9]), .B2(EX__n1256), .Y(EX__n1543) );
  INVx1_ASAP7_75t_R EX___U1245 ( .A(EX__n685), .Y(EX__n952) );
  BUFx10_ASAP7_75t_R EX___U1246 ( .A(EX__n954), .Y(EX__n953) );
  BUFx4f_ASAP7_75t_R EX___U1247 ( .A(EX__n648), .Y(EX__n954) );
  BUFx16f_ASAP7_75t_R EX___U1248 ( .A(EX__n650), .Y(EX__n1211) );
  BUFx2_ASAP7_75t_R EX___U1249 ( .A(EX__n1213), .Y(EX__n956) );
  BUFx10_ASAP7_75t_R EX___U1250 ( .A(EX__n958), .Y(EX__n957) );
  BUFx4f_ASAP7_75t_R EX___U1251 ( .A(EX__n465), .Y(EX__n958) );
  BUFx2_ASAP7_75t_R EX___U1252 ( .A(EX__n1168), .Y(EX__n959) );
  BUFx3_ASAP7_75t_R EX___U1253 ( .A(ID_EX_imm[30]), .Y(EX__n1475) );
  OR2x2_ASAP7_75t_R EX___U1254 ( .A(EX__n1336), .B(EX__n1464), .Y(EX__n1466) );
  INVx2_ASAP7_75t_R EX___U1255 ( .A(EX__n447), .Y(EX__n961) );
  OA22x2_ASAP7_75t_R EX___U1256 ( .A1(EX__n1365), .A2(EX__n454), .B1(EX__n1611), .B2(EX__n1350), 
        .Y(EX__n1465) );
  INVx2_ASAP7_75t_R EX___U1257 ( .A(EX__n449), .Y(EX__n962) );
  CKINVDCx20_ASAP7_75t_R EX___U1258 ( .A(EX__n292), .Y(EX__n963) );
  CKINVDCx20_ASAP7_75t_R EX___U1259 ( .A(EX__n963), .Y(EX__n964) );
  OR2x2_ASAP7_75t_R EX___U1260 ( .A(EX__n1329), .B(EX__n1422), .Y(EX__n1424) );
  INVx2_ASAP7_75t_R EX___U1261 ( .A(EX__n163), .Y(EX__n966) );
  OA22x2_ASAP7_75t_R EX___U1262 ( .A1(EX__n1361), .A2(EX__n784), .B1(EX__n1597), .B2(EX__n1348), 
        .Y(EX__n1423) );
  INVx2_ASAP7_75t_R EX___U1263 ( .A(EX__n165), .Y(EX__n967) );
  CKINVDCx20_ASAP7_75t_R EX___U1264 ( .A(EX__n98), .Y(EX__n968) );
  CKINVDCx20_ASAP7_75t_R EX___U1265 ( .A(EX__n968), .Y(EX__n969) );
  OR2x2_ASAP7_75t_R EX___U1266 ( .A(EX__n1333), .B(EX__n1446), .Y(EX__n1448) );
  INVx2_ASAP7_75t_R EX___U1267 ( .A(EX__n212), .Y(EX__n971) );
  OA22x2_ASAP7_75t_R EX___U1268 ( .A1(EX__n1364), .A2(EX__n511), .B1(EX__n1605), .B2(EX__n458), .Y(
        n1447) );
  INVx2_ASAP7_75t_R EX___U1269 ( .A(EX__n214), .Y(EX__n972) );
  CKINVDCx20_ASAP7_75t_R EX___U1270 ( .A(EX__n217), .Y(EX__n973) );
  BUFx4f_ASAP7_75t_R EX___U1271 ( .A(ID_EX_imm[16]), .Y(EX__n1523) );
  INVx2_ASAP7_75t_R EX___U1272 ( .A(EX__n1523), .Y(EX__n975) );
  OA22x2_ASAP7_75t_R EX___U1273 ( .A1(EX__n976), .A2(EX__n1311), .B1(EX__n73), .B2(EX__n975), .Y(
        input_data_2[16]) );
  OA22x2_ASAP7_75t_R EX___U1274 ( .A1(EX__n979), .A2(EX__n407), .B1(EX__n1295), .B2(EX__n1489), .Y(
        input_data_2[26]) );
  INVx1_ASAP7_75t_R EX___U1275 ( .A(EX__n1490), .Y(EX__n979) );
  INVx1_ASAP7_75t_R EX___U1276 ( .A(EX__n1045), .Y(EX__n980) );
  BUFx3_ASAP7_75t_R EX___U1277 ( .A(EX__n988), .Y(EX__n987) );
  BUFx2_ASAP7_75t_R EX___U1278 ( .A(EX__n1513), .Y(EX__n988) );
  INVx1_ASAP7_75t_R EX___U1279 ( .A(EX__n868), .Y(EX__n991) );
  BUFx3_ASAP7_75t_R EX___U1280 ( .A(forwarding_MEM_WB[0]), .Y(EX__n1574) );
  INVx1_ASAP7_75t_R EX___U1281 ( .A(EX__n870), .Y(EX__n992) );
  BUFx3_ASAP7_75t_R EX___U1282 ( .A(forwarding_MEM_WB[21]), .Y(EX__n1506) );
  BUFx3_ASAP7_75t_R EX___U1283 ( .A(forwarding_MEM_WB[8]), .Y(EX__n1547) );
  INVx1_ASAP7_75t_R EX___U1284 ( .A(EX__n875), .Y(EX__n996) );
  INVx1_ASAP7_75t_R EX___U1285 ( .A(EX__n873), .Y(EX__n998) );
  BUFx3_ASAP7_75t_R EX___U1286 ( .A(EX__n807), .Y(EX__n1000) );
  OA21x2_ASAP7_75t_R EX___U1287 ( .A1(EX__n627), .A2(EX__n35), .B(EX__n1002), .Y(EX__n1638) );
  INVx2_ASAP7_75t_R EX___U1288 ( .A(EX__n414), .Y(EX_read_reg_data_2[4]) );
  AO22x2_ASAP7_75t_R EX___U1289 ( .A1(forwarding_EX_MEM[4]), .A2(EX__n1274), .B1(
        ID_EX_read_reg_data_2[4]), .B2(EX__n344), .Y(EX__n1562) );
  INVx1_ASAP7_75t_R EX___U1290 ( .A(EX__n416), .Y(EX__n1002) );
  AO22x2_ASAP7_75t_R EX___U1291 ( .A1(forwarding_EX_MEM[27]), .A2(EX__n1266), .B1(
        ID_EX_read_reg_data_2[27]), .B2(EX__n761), .Y(EX__n1484) );
  OA21x2_ASAP7_75t_R EX___U1292 ( .A1(EX__n1286), .A2(EX__n1191), .B(EX__n1005), .Y(EX__n1620) );
  AO22x2_ASAP7_75t_R EX___U1293 ( .A1(forwarding_EX_MEM[23]), .A2(EX__n1267), .B1(
        ID_EX_read_reg_data_2[23]), .B2(EX__n1260), .Y(EX__n1498) );
  INVx1_ASAP7_75t_R EX___U1294 ( .A(EX__n570), .Y(EX__n1005) );
  AO22x2_ASAP7_75t_R EX___U1295 ( .A1(forwarding_EX_MEM[6]), .A2(EX__n1273), .B1(
        ID_EX_read_reg_data_2[6]), .B2(EX__n295), .Y(EX__n1554) );
  INVx1_ASAP7_75t_R EX___U1296 ( .A(EX__n727), .Y(EX__n1006) );
  OR2x2_ASAP7_75t_R EX___U1297 ( .A(EX__n1322), .B(EX__n1374), .Y(EX__n1376) );
  INVx2_ASAP7_75t_R EX___U1298 ( .A(EX__n594), .Y(EX__n1007) );
  OA22x2_ASAP7_75t_R EX___U1299 ( .A1(EX__n1041), .A2(EX__n84), .B1(EX__n1581), .B2(EX__n264), .Y(
        n1375) );
  INVx2_ASAP7_75t_R EX___U1300 ( .A(EX__n596), .Y(EX__n1008) );
  CKINVDCx20_ASAP7_75t_R EX___U1301 ( .A(EX__n370), .Y(EX__n1009) );
  CKINVDCx20_ASAP7_75t_R EX___U1302 ( .A(EX__n1009), .Y(EX__n1010) );
  OR2x2_ASAP7_75t_R EX___U1303 ( .A(EX__n1336), .B(EX__n1461), .Y(EX__n1463) );
  INVx2_ASAP7_75t_R EX___U1304 ( .A(EX__n372), .Y(EX__n1012) );
  OA22x2_ASAP7_75t_R EX___U1305 ( .A1(EX__n1365), .A2(EX__n769), .B1(EX__n1610), .B2(EX__n1350), 
        .Y(EX__n1462) );
  INVx2_ASAP7_75t_R EX___U1306 ( .A(EX__n374), .Y(EX__n1013) );
  CKINVDCx20_ASAP7_75t_R EX___U1307 ( .A(EX__n209), .Y(EX__n1014) );
  CKINVDCx20_ASAP7_75t_R EX___U1308 ( .A(EX__n1014), .Y(EX__n1015) );
  OR2x2_ASAP7_75t_R EX___U1309 ( .A(EX__n1330), .B(EX__n1425), .Y(EX__n1427) );
  INVx2_ASAP7_75t_R EX___U1310 ( .A(EX__n184), .Y(EX__n1017) );
  OA22x2_ASAP7_75t_R EX___U1311 ( .A1(EX__n1362), .A2(EX__n943), .B1(EX__n1598), .B2(EX__n255), .Y(
        n1426) );
  INVx2_ASAP7_75t_R EX___U1312 ( .A(EX__n186), .Y(EX__n1018) );
  CKINVDCx20_ASAP7_75t_R EX___U1313 ( .A(EX__n112), .Y(EX__n1019) );
  CKINVDCx20_ASAP7_75t_R EX___U1314 ( .A(EX__n1019), .Y(EX__n1020) );
  OR2x2_ASAP7_75t_R EX___U1315 ( .A(EX__n1325), .B(EX__n1398), .Y(EX__n1400) );
  INVx2_ASAP7_75t_R EX___U1316 ( .A(EX__n354), .Y(EX__n1022) );
  OA22x2_ASAP7_75t_R EX___U1317 ( .A1(EX__n1359), .A2(EX__n702), .B1(EX__n1132), .B2(EX__n1346), 
        .Y(EX__n1399) );
  INVx2_ASAP7_75t_R EX___U1318 ( .A(EX__n356), .Y(EX__n1023) );
  CKINVDCx20_ASAP7_75t_R EX___U1319 ( .A(EX__n359), .Y(EX__n1024) );
  OR2x2_ASAP7_75t_R EX___U1320 ( .A(EX__n1332), .B(EX__n1437), .Y(EX__n1439) );
  INVx2_ASAP7_75t_R EX___U1321 ( .A(EX__n540), .Y(EX__n1026) );
  OA22x2_ASAP7_75t_R EX___U1322 ( .A1(EX__n1363), .A2(EX__n1040), .B1(EX__n1602), .B2(EX__n257), 
        .Y(EX__n1438) );
  INVx2_ASAP7_75t_R EX___U1323 ( .A(EX__n542), .Y(EX__n1027) );
  CKINVDCx20_ASAP7_75t_R EX___U1324 ( .A(EX__n141), .Y(EX__n1028) );
  CKINVDCx20_ASAP7_75t_R EX___U1325 ( .A(EX__n1028), .Y(EX__n1029) );
  OA22x2_ASAP7_75t_R EX___U1326 ( .A1(EX__n1032), .A2(EX__n1311), .B1(EX__n1297), .B2(EX__n1511), 
        .Y(input_data_2[20]) );
  INVx1_ASAP7_75t_R EX___U1327 ( .A(EX__n1512), .Y(EX__n1032) );
  OA22x2_ASAP7_75t_R EX___U1328 ( .A1(EX__n1034), .A2(EX__n1321), .B1(EX__n1295), .B2(EX__n1482), 
        .Y(input_data_2[28]) );
  INVx1_ASAP7_75t_R EX___U1329 ( .A(EX__n1483), .Y(EX__n1034) );
  BUFx4f_ASAP7_75t_R EX___U1330 ( .A(EX__n1488), .Y(EX__n1036) );
  INVx1_ASAP7_75t_R EX___U1331 ( .A(ID_EX_read_reg_data_1[23]), .Y(EX__n1588) );
  INVx1_ASAP7_75t_R EX___U1332 ( .A(EX__n866), .Y(EX__n1041) );
  BUFx3_ASAP7_75t_R EX___U1333 ( .A(forwarding_MEM_WB[17]), .Y(EX__n1519) );
  INVx1_ASAP7_75t_R EX___U1334 ( .A(EX__n981), .Y(EX__n1044) );
  AO22x2_ASAP7_75t_R EX___U1335 ( .A1(forwarding_EX_MEM[25]), .A2(EX__n1267), .B1(
        ID_EX_read_reg_data_2[25]), .B2(EX__n1258), .Y(EX__n1491) );
  OA21x2_ASAP7_75t_R EX___U1336 ( .A1(EX__n1284), .A2(EX__n26), .B(EX__n1049), .Y(EX__n1628) );
  AO22x2_ASAP7_75t_R EX___U1337 ( .A1(forwarding_EX_MEM[15]), .A2(EX__n1270), .B1(
        ID_EX_read_reg_data_2[15]), .B2(EX__n1255), .Y(EX__n1524) );
  INVx1_ASAP7_75t_R EX___U1338 ( .A(EX__n642), .Y(EX__n1049) );
  AO22x2_ASAP7_75t_R EX___U1339 ( .A1(forwarding_EX_MEM[22]), .A2(EX__n1268), .B1(
        ID_EX_read_reg_data_2[22]), .B2(EX__n325), .Y(EX__n1501) );
  INVx2_ASAP7_75t_R EX___U1340 ( .A(EX__n644), .Y(EX_read_reg_data_2[13]) );
  AO22x2_ASAP7_75t_R EX___U1341 ( .A1(forwarding_EX_MEM[13]), .A2(EX__n1271), .B1(
        ID_EX_read_reg_data_2[13]), .B2(EX__n1259), .Y(EX__n1531) );
  OA21x2_ASAP7_75t_R EX___U1342 ( .A1(EX__n1282), .A2(EX__n61), .B(EX__n1053), .Y(EX__n1636) );
  AO22x2_ASAP7_75t_R EX___U1343 ( .A1(forwarding_EX_MEM[7]), .A2(EX__n1273), .B1(
        ID_EX_read_reg_data_2[7]), .B2(EX__n630), .Y(EX__n1550) );
  INVx1_ASAP7_75t_R EX___U1344 ( .A(EX__n657), .Y(EX__n1053) );
  BUFx10_ASAP7_75t_R EX___U1345 ( .A(EX__n1055), .Y(EX__n1054) );
  BUFx4f_ASAP7_75t_R EX___U1346 ( .A(EX__n713), .Y(EX__n1055) );
  BUFx16f_ASAP7_75t_R EX___U1347 ( .A(EX__n715), .Y(EX__n1125) );
  CKINVDCx20_ASAP7_75t_R EX___U1348 ( .A(EX__n1125), .Y(EX__n1056) );
  BUFx2_ASAP7_75t_R EX___U1349 ( .A(EX__n1126), .Y(EX__n1057) );
  OR2x2_ASAP7_75t_R EX___U1350 ( .A(EX__n1335), .B(EX__n1455), .Y(EX__n1457) );
  INVx2_ASAP7_75t_R EX___U1351 ( .A(EX__n236), .Y(EX__n1058) );
  OA22x2_ASAP7_75t_R EX___U1352 ( .A1(EX__n991), .A2(EX__n267), .B1(EX__n1608), .B2(EX__n1348), .Y(
        n1456) );
  INVx2_ASAP7_75t_R EX___U1353 ( .A(EX__n238), .Y(EX__n1059) );
  CKINVDCx20_ASAP7_75t_R EX___U1354 ( .A(EX__n241), .Y(EX__n1060) );
  OR2x2_ASAP7_75t_R EX___U1355 ( .A(EX__n1324), .B(EX__n1392), .Y(EX__n1394) );
  INVx2_ASAP7_75t_R EX___U1356 ( .A(EX__n377), .Y(EX__n1062) );
  OA22x2_ASAP7_75t_R EX___U1357 ( .A1(EX__n1358), .A2(EX__n1133), .B1(EX__n1587), .B2(EX__n1345), 
        .Y(EX__n1393) );
  INVx2_ASAP7_75t_R EX___U1358 ( .A(EX__n379), .Y(EX__n1063) );
  CKINVDCx20_ASAP7_75t_R EX___U1359 ( .A(EX__n382), .Y(EX__n1064) );
  OR2x2_ASAP7_75t_R EX___U1360 ( .A(EX__n1326), .B(EX__n1404), .Y(EX__n1406) );
  INVx2_ASAP7_75t_R EX___U1361 ( .A(EX__n156), .Y(EX__n1066) );
  OA22x2_ASAP7_75t_R EX___U1362 ( .A1(EX__n1359), .A2(EX__n479), .B1(EX__n1591), .B2(EX__n1346), 
        .Y(EX__n1405) );
  INVx2_ASAP7_75t_R EX___U1363 ( .A(EX__n158), .Y(EX__n1067) );
  CKINVDCx20_ASAP7_75t_R EX___U1364 ( .A(EX__n161), .Y(EX__n1068) );
  OR2x2_ASAP7_75t_R EX___U1365 ( .A(EX__n1328), .B(EX__n1416), .Y(EX__n1418) );
  INVx2_ASAP7_75t_R EX___U1366 ( .A(EX__n327), .Y(EX__n1070) );
  OA22x2_ASAP7_75t_R EX___U1367 ( .A1(EX__n1361), .A2(EX__n733), .B1(EX__n1595), .B2(EX__n1348), 
        .Y(EX__n1417) );
  INVx2_ASAP7_75t_R EX___U1368 ( .A(EX__n329), .Y(EX__n1071) );
  CKINVDCx20_ASAP7_75t_R EX___U1369 ( .A(EX__n259), .Y(EX__n1072) );
  CKINVDCx20_ASAP7_75t_R EX___U1370 ( .A(EX__n1072), .Y(EX__n1073) );
  OA22x2_ASAP7_75t_R EX___U1371 ( .A1(EX__n1076), .A2(EX__n1311), .B1(EX__n1507), .B2(EX__n1297), 
        .Y(input_data_2[21]) );
  INVx1_ASAP7_75t_R EX___U1372 ( .A(EX__n1508), .Y(EX__n1076) );
  OA22x2_ASAP7_75t_R EX___U1373 ( .A1(EX__n620), .A2(EX__n1314), .B1(EX__n1301), .B2(EX__n1078), 
        .Y(input_data_2[8]) );
  BUFx2_ASAP7_75t_R EX___U1374 ( .A(EX__n1548), .Y(EX__n1078) );
  BUFx2_ASAP7_75t_R EX___U1375 ( .A(EX_read_reg_data_2[8]), .Y(EX__n1549) );
  INVx1_ASAP7_75t_R EX___U1376 ( .A(EX__n1549), .Y(EX__n1079) );
  BUFx2_ASAP7_75t_R EX___U1377 ( .A(ID_EX_read_reg_data_1[5]), .Y(EX__n1606) );
  INVx1_ASAP7_75t_R EX___U1378 ( .A(EX__n1606), .Y(EX__n1080) );
  BUFx2_ASAP7_75t_R EX___U1379 ( .A(ID_EX_read_reg_data_1[25]), .Y(EX__n1586) );
  INVx1_ASAP7_75t_R EX___U1380 ( .A(EX__n1586), .Y(EX__n1081) );
  BUFx12f_ASAP7_75t_R EX___U1381 ( .A(EX__n1257), .Y(EX__n1262) );
  BUFx12f_ASAP7_75t_R EX___U1382 ( .A(EX__n1264), .Y(EX__n1263) );
  BUFx12f_ASAP7_75t_R EX___U1383 ( .A(EX__n485), .Y(EX__n1280) );
  INVx3_ASAP7_75t_R EX___U1384 ( .A(ForwardA[1]), .Y(EX__n1578) );
  BUFx12f_ASAP7_75t_R EX___U1385 ( .A(EX__n482), .Y(EX__n1085) );
  AND2x2_ASAP7_75t_R EX___U1386 ( .A(ForwardB[0]), .B(EX__n1467), .Y(EX__n1575) );
  INVx2_ASAP7_75t_R EX___U1387 ( .A(EX__n483), .Y(EX__n1086) );
  BUFx12f_ASAP7_75t_R EX___U1388 ( .A(EX__n760), .Y(EX__n1293) );
  BUFx8_ASAP7_75t_R EX___U1389 ( .A(EX__n1086), .Y(EX__n1294) );
  CKINVDCx5p33_ASAP7_75t_R EX___U1390 ( .A(EX__n1332), .Y(EX__n1087) );
  INVx2_ASAP7_75t_R EX___U1391 ( .A(EX__n1087), .Y(EX__n1334) );
  INVx3_ASAP7_75t_R EX___U1392 ( .A(EX__n1087), .Y(EX__n1333) );
  BUFx12f_ASAP7_75t_R EX___U1393 ( .A(EX__n253), .Y(EX__n1337) );
  OR2x2_ASAP7_75t_R EX___U1394 ( .A(EX__n1322), .B(EX__n1371), .Y(EX__n1373) );
  INVx2_ASAP7_75t_R EX___U1395 ( .A(EX__n504), .Y(EX__n1088) );
  OA22x2_ASAP7_75t_R EX___U1396 ( .A1(EX__n85), .A2(EX__n436), .B1(EX__n1580), .B2(EX__n265), .Y(
        n1372) );
  INVx2_ASAP7_75t_R EX___U1397 ( .A(EX__n506), .Y(EX__n1089) );
  CKINVDCx20_ASAP7_75t_R EX___U1398 ( .A(EX__n409), .Y(EX__n1090) );
  CKINVDCx20_ASAP7_75t_R EX___U1399 ( .A(EX__n1090), .Y(EX__n1091) );
  OR2x2_ASAP7_75t_R EX___U1400 ( .A(EX__n1335), .B(EX__n1458), .Y(EX__n1460) );
  INVx2_ASAP7_75t_R EX___U1401 ( .A(EX__n740), .Y(EX__n1093) );
  OA22x2_ASAP7_75t_R EX___U1402 ( .A1(EX__n1364), .A2(EX__n768), .B1(EX__n1609), .B2(EX__n289), .Y(
        n1459) );
  INVx2_ASAP7_75t_R EX___U1403 ( .A(EX__n742), .Y(EX__n1094) );
  OR2x2_ASAP7_75t_R EX___U1404 ( .A(EX__n1323), .B(EX__n1386), .Y(EX__n1388) );
  INVx2_ASAP7_75t_R EX___U1405 ( .A(EX__n496), .Y(EX__n1098) );
  OA22x2_ASAP7_75t_R EX___U1406 ( .A1(EX__n1190), .A2(EX__n1357), .B1(EX__n1585), .B2(EX__n459), 
        .Y(EX__n1387) );
  INVx2_ASAP7_75t_R EX___U1407 ( .A(EX__n498), .Y(EX__n1099) );
  CKINVDCx20_ASAP7_75t_R EX___U1408 ( .A(EX__n501), .Y(EX__n1100) );
  OR2x2_ASAP7_75t_R EX___U1409 ( .A(EX__n1327), .B(EX__n1407), .Y(EX__n1409) );
  INVx2_ASAP7_75t_R EX___U1410 ( .A(EX__n745), .Y(EX__n1102) );
  OA22x2_ASAP7_75t_R EX___U1411 ( .A1(EX__n1135), .A2(EX__n1360), .B1(EX__n1592), .B2(EX__n1347), 
        .Y(EX__n1408) );
  INVx2_ASAP7_75t_R EX___U1412 ( .A(EX__n747), .Y(EX__n1103) );
  CKINVDCx20_ASAP7_75t_R EX___U1413 ( .A(EX__n609), .Y(EX__n1104) );
  OR2x2_ASAP7_75t_R EX___U1414 ( .A(EX__n1330), .B(EX__n1428), .Y(EX__n1430) );
  INVx2_ASAP7_75t_R EX___U1415 ( .A(EX__n300), .Y(EX__n1107) );
  OA22x2_ASAP7_75t_R EX___U1416 ( .A1(EX__n1362), .A2(EX__n803), .B1(EX__n1599), .B2(EX__n263), .Y(
        n1429) );
  INVx2_ASAP7_75t_R EX___U1417 ( .A(EX__n302), .Y(EX__n1108) );
  CKINVDCx20_ASAP7_75t_R EX___U1418 ( .A(EX__n234), .Y(EX__n1109) );
  OR2x2_ASAP7_75t_R EX___U1419 ( .A(EX__n1333), .B(EX__n1443), .Y(EX__n1445) );
  INVx2_ASAP7_75t_R EX___U1420 ( .A(EX__n771), .Y(EX__n1111) );
  OA22x2_ASAP7_75t_R EX___U1421 ( .A1(EX__n1364), .A2(EX__n604), .B1(EX__n1604), .B2(EX__n1348), 
        .Y(EX__n1444) );
  INVx2_ASAP7_75t_R EX___U1422 ( .A(EX__n773), .Y(EX__n1112) );
  CKINVDCx20_ASAP7_75t_R EX___U1423 ( .A(EX__n1115), .Y(EX__n1113) );
  CKINVDCx20_ASAP7_75t_R EX___U1424 ( .A(EX__n588), .Y(EX__n1114) );
  BUFx16f_ASAP7_75t_R EX___U1425 ( .A(EX__n770), .Y(EX__n1115) );
  INVx2_ASAP7_75t_R EX___U1426 ( .A(EX__n1532), .Y(EX__n1116) );
  BUFx2_ASAP7_75t_R EX___U1427 ( .A(EX_read_reg_data_2[13]), .Y(EX__n1533) );
  OA22x2_ASAP7_75t_R EX___U1428 ( .A1(EX__n764), .A2(EX__n1313), .B1(EX__n1300), .B2(EX__n1116), 
        .Y(input_data_2[13]) );
  INVx2_ASAP7_75t_R EX___U1429 ( .A(EX__n1570), .Y(EX__n1119) );
  BUFx4f_ASAP7_75t_R EX___U1430 ( .A(EX__n695), .Y(EX__n1571) );
  INVx2_ASAP7_75t_R EX___U1431 ( .A(EX__n1571), .Y(EX__n1120) );
  OA22x2_ASAP7_75t_R EX___U1432 ( .A1(EX__n1120), .A2(EX__n1315), .B1(EX__n1303), .B2(EX__n1119), 
        .Y(input_data_2[1]) );
  OA22x2_ASAP7_75t_R EX___U1433 ( .A1(EX__n1124), .A2(EX__n1309), .B1(EX__n363), .B2(EX__n1478), 
        .Y(input_data_2[29]) );
  INVx2_ASAP7_75t_R EX___U1434 ( .A(ID_EX_imm[29]), .Y(EX__n1478) );
  OA22x2_ASAP7_75t_R EX___U1435 ( .A1(EX__n1057), .A2(EX__n1310), .B1(EX__n1499), .B2(EX__n1296), 
        .Y(input_data_2[23]) );
  OA22x2_ASAP7_75t_R EX___U1436 ( .A1(EX__n791), .A2(EX__n1312), .B1(EX__n1298), .B2(EX__n1128), 
        .Y(input_data_2[17]) );
  INVx1_ASAP7_75t_R EX___U1437 ( .A(EX__n1520), .Y(EX__n1128) );
  INVx1_ASAP7_75t_R EX___U1438 ( .A(EX__n1521), .Y(EX__n1129) );
  OA22x2_ASAP7_75t_R EX___U1439 ( .A1(EX__n799), .A2(EX__n1312), .B1(EX__n1560), .B2(EX__n1302), 
        .Y(input_data_2[5]) );
  BUFx2_ASAP7_75t_R EX___U1440 ( .A(ID_EX_read_reg_data_1[22]), .Y(EX__n1589) );
  INVx1_ASAP7_75t_R EX___U1441 ( .A(EX__n1589), .Y(EX__n1132) );
  INVx1_ASAP7_75t_R EX___U1442 ( .A(EX__n1038), .Y(EX__n1135) );
  OA21x2_ASAP7_75t_R EX___U1443 ( .A1(EX__n1288), .A2(EX__n785), .B(EX__n1137), .Y(EX__n1612) );
  INVx2_ASAP7_75t_R EX___U1444 ( .A(EX__n705), .Y(EX_read_reg_data_2[31]) );
  AO22x2_ASAP7_75t_R EX___U1445 ( .A1(forwarding_EX_MEM[31]), .A2(EX__n1265), .B1(
        ID_EX_read_reg_data_2[31]), .B2(EX__n1255), .Y(EX__n1470) );
  INVx1_ASAP7_75t_R EX___U1446 ( .A(EX__n707), .Y(EX__n1137) );
  INVx2_ASAP7_75t_R EX___U1447 ( .A(EX__n830), .Y(EX_read_reg_data_2[26]) );
  AO22x2_ASAP7_75t_R EX___U1448 ( .A1(forwarding_EX_MEM[26]), .A2(EX__n1266), .B1(
        ID_EX_read_reg_data_2[26]), .B2(EX__n631), .Y(EX__n1487) );
  OA21x2_ASAP7_75t_R EX___U1449 ( .A1(EX__n1286), .A2(EX__n30), .B(EX__n1140), .Y(EX__n1622) );
  AO22x2_ASAP7_75t_R EX___U1450 ( .A1(forwarding_EX_MEM[21]), .A2(EX__n1268), .B1(
        ID_EX_read_reg_data_2[21]), .B2(EX__n291), .Y(EX__n1505) );
  INVx1_ASAP7_75t_R EX___U1451 ( .A(EX__n906), .Y(EX__n1140) );
  INVx2_ASAP7_75t_R EX___U1452 ( .A(EX__n532), .Y(EX_read_reg_data_2[8]) );
  AO22x2_ASAP7_75t_R EX___U1453 ( .A1(forwarding_EX_MEM[8]), .A2(EX__n1272), .B1(
        ID_EX_read_reg_data_2[8]), .B2(EX__n1256), .Y(EX__n1546) );
  OA21x2_ASAP7_75t_R EX___U1454 ( .A1(EX__n1292), .A2(EX__n863), .B(EX__n1143), .Y(EX__n1637) );
  AO22x2_ASAP7_75t_R EX___U1455 ( .A1(forwarding_EX_MEM[5]), .A2(EX__n1273), .B1(
        ID_EX_read_reg_data_2[5]), .B2(EX__n1256), .Y(EX__n1558) );
  INVx1_ASAP7_75t_R EX___U1456 ( .A(EX__n941), .Y(EX__n1143) );
  OA21x2_ASAP7_75t_R EX___U1457 ( .A1(EX__n1284), .A2(EX__n1043), .B(EX__n1145), .Y(EX__n1626) );
  INVx2_ASAP7_75t_R EX___U1458 ( .A(EX__n931), .Y(EX_read_reg_data_2[17]) );
  AO22x2_ASAP7_75t_R EX___U1459 ( .A1(forwarding_EX_MEM[17]), .A2(EX__n1269), .B1(
        ID_EX_read_reg_data_2[17]), .B2(EX__n1255), .Y(EX__n1518) );
  INVx1_ASAP7_75t_R EX___U1460 ( .A(EX__n933), .Y(EX__n1145) );
  OA21x2_ASAP7_75t_R EX___U1461 ( .A1(EX__n1283), .A2(EX__n33), .B(EX__n1147), .Y(EX__n1631) );
  AO22x2_ASAP7_75t_R EX___U1462 ( .A1(forwarding_EX_MEM[12]), .A2(EX__n1271), .B1(
        ID_EX_read_reg_data_2[12]), .B2(EX__n1264), .Y(EX__n1534) );
  INVx1_ASAP7_75t_R EX___U1463 ( .A(EX__n937), .Y(EX__n1147) );
  OR2x6_ASAP7_75t_R EX___U1464 ( .A(EX__n1062), .B(EX__n1063), .Y(input_A[24]) );
  OR2x6_ASAP7_75t_R EX___U1465 ( .A(EX__n1022), .B(EX__n1023), .Y(input_A[22]) );
  OR2x6_ASAP7_75t_R EX___U1466 ( .A(EX__n1102), .B(EX__n1103), .Y(input_A[19]) );
  XOR2x2_ASAP7_75t_R EX___U1467 ( .A(ForwardA[0]), .B(ForwardA[1]), .Y(EX__n139) );
  BUFx2_ASAP7_75t_R EX___U1468 ( .A(EX__n5), .Y(EX__n1148) );
  OR2x2_ASAP7_75t_R EX___U1469 ( .A(EX__n1331), .B(EX__n1431), .Y(EX__n1433) );
  INVx2_ASAP7_75t_R EX___U1470 ( .A(EX__n844), .Y(EX__n1149) );
  OA22x2_ASAP7_75t_R EX___U1471 ( .A1(EX__n1362), .A2(EX__n783), .B1(EX__n1189), .B2(EX__n288), .Y(
        n1432) );
  INVx2_ASAP7_75t_R EX___U1472 ( .A(EX__n846), .Y(EX__n1150) );
  CKINVDCx20_ASAP7_75t_R EX___U1473 ( .A(EX__n1153), .Y(EX__n1151) );
  CKINVDCx20_ASAP7_75t_R EX___U1474 ( .A(EX__n494), .Y(EX__n1152) );
  BUFx16f_ASAP7_75t_R EX___U1475 ( .A(EX__n843), .Y(EX__n1153) );
  INVx2_ASAP7_75t_R EX___U1476 ( .A(EX__n983), .Y(EX__n1154) );
  INVx2_ASAP7_75t_R EX___U1477 ( .A(EX__n1493), .Y(EX__n1155) );
  OA22x2_ASAP7_75t_R EX___U1478 ( .A1(EX__n1154), .A2(EX__n1310), .B1(EX__n1296), .B2(EX__n1155), 
        .Y(input_data_2[25]) );
  OR2x2_ASAP7_75t_R EX___U1479 ( .A(EX__n1323), .B(EX__n1383), .Y(EX__n1385) );
  INVx2_ASAP7_75t_R EX___U1480 ( .A(EX__n278), .Y(EX__n1158) );
  OA22x2_ASAP7_75t_R EX___U1481 ( .A1(EX__n1357), .A2(EX__n510), .B1(EX__n1584), .B2(EX__n1353), 
        .Y(EX__n1384) );
  INVx2_ASAP7_75t_R EX___U1482 ( .A(EX__n280), .Y(EX__n1159) );
  CKINVDCx20_ASAP7_75t_R EX___U1483 ( .A(EX__n283), .Y(EX__n1160) );
  OA22x2_ASAP7_75t_R EX___U1484 ( .A1(EX__n738), .A2(EX__n1311), .B1(EX__n1503), .B2(EX__n1297), 
        .Y(input_data_2[22]) );
  OA22x2_ASAP7_75t_R EX___U1485 ( .A1(EX__n1166), .A2(EX__n1314), .B1(EX__n1301), .B2(EX__n1165), 
        .Y(input_data_2[10]) );
  INVx1_ASAP7_75t_R EX___U1486 ( .A(EX__n1541), .Y(EX__n1165) );
  INVx1_ASAP7_75t_R EX___U1487 ( .A(EX__n1542), .Y(EX__n1166) );
  OA22x2_ASAP7_75t_R EX___U1488 ( .A1(EX__n959), .A2(EX__n1309), .B1(EX__n1308), .B2(EX__n1169), 
        .Y(input_data_2[30]) );
  INVx1_ASAP7_75t_R EX___U1489 ( .A(EX__n1475), .Y(EX__n1169) );
  OA22x2_ASAP7_75t_R EX___U1490 ( .A1(EX__n795), .A2(EX__n1309), .B1(EX__n74), .B2(EX__n1171), .Y(
        input_data_2[14]) );
  INVx1_ASAP7_75t_R EX___U1491 ( .A(EX__n1529), .Y(EX__n1171) );
  CKINVDCx20_ASAP7_75t_R EX___U1492 ( .A(EX__n428), .Y(EX__n1173) );
  CKINVDCx20_ASAP7_75t_R EX___U1493 ( .A(EX__n600), .Y(EX__n1174) );
  OR2x2_ASAP7_75t_R EX___U1494 ( .A(EX__n1334), .B(EX__n1452), .Y(EX__n1454) );
  INVx1_ASAP7_75t_R EX___U1495 ( .A(EX__n601), .Y(EX__n1176) );
  OA22x2_ASAP7_75t_R EX___U1496 ( .A1(EX__n1358), .A2(EX__n528), .B1(EX__n1607), .B2(EX__n1351), 
        .Y(EX__n1453) );
  INVx1_ASAP7_75t_R EX___U1497 ( .A(EX__n602), .Y(EX__n1177) );
  OR2x4_ASAP7_75t_R EX___U1498 ( .A(EX__n1176), .B(EX__n1177), .Y(input_A[4]) );
  CKINVDCx20_ASAP7_75t_R EX___U1499 ( .A(EX__n663), .Y(EX__n1178) );
  OR2x2_ASAP7_75t_R EX___U1500 ( .A(EX__n1325), .B(EX__n1395), .Y(EX__n1397) );
  INVx1_ASAP7_75t_R EX___U1501 ( .A(EX__n664), .Y(EX__n1180) );
  OA22x2_ASAP7_75t_R EX___U1502 ( .A1(EX__n1358), .A2(EX__n881), .B1(EX__n1588), .B2(EX__n1345), 
        .Y(EX__n1396) );
  INVx1_ASAP7_75t_R EX___U1503 ( .A(EX__n665), .Y(EX__n1181) );
  OR2x4_ASAP7_75t_R EX___U1504 ( .A(EX__n1180), .B(EX__n1181), .Y(input_A[23]) );
  CKINVDCx20_ASAP7_75t_R EX___U1505 ( .A(EX__n366), .Y(EX__n1182) );
  OR2x2_ASAP7_75t_R EX___U1506 ( .A(EX__n1327), .B(EX__n1410), .Y(EX__n1412) );
  INVx1_ASAP7_75t_R EX___U1507 ( .A(EX__n367), .Y(EX__n1184) );
  OA22x2_ASAP7_75t_R EX___U1508 ( .A1(EX__n1360), .A2(EX__n882), .B1(EX__n1593), .B2(EX__n1347), 
        .Y(EX__n1411) );
  INVx1_ASAP7_75t_R EX___U1509 ( .A(EX__n368), .Y(EX__n1185) );
  OR2x4_ASAP7_75t_R EX___U1510 ( .A(EX__n1184), .B(EX__n1185), .Y(input_A[18]) );
  OA22x2_ASAP7_75t_R EX___U1511 ( .A1(EX__n896), .A2(EX__n1315), .B1(EX__n1303), .B2(EX__n1187), 
        .Y(input_data_2[0]) );
  INVx1_ASAP7_75t_R EX___U1512 ( .A(EX__n1576), .Y(EX__n1187) );
  INVx1_ASAP7_75t_R EX___U1513 ( .A(EX__n1577), .Y(EX__n1188) );
  BUFx2_ASAP7_75t_R EX___U1514 ( .A(ID_EX_read_reg_data_1[11]), .Y(EX__n1600) );
  INVx1_ASAP7_75t_R EX___U1515 ( .A(EX__n1600), .Y(EX__n1189) );
  OR2x6_ASAP7_75t_R EX___U1516 ( .A(EX__n1088), .B(EX__n1089), .Y(input_A[31]) );
  BUFx3_ASAP7_75t_R EX___U1517 ( .A(forwarding_MEM_WB[26]), .Y(EX__n1488) );
  INVx1_ASAP7_75t_R EX___U1518 ( .A(EX__n1035), .Y(EX__n1190) );
  INVx2_ASAP7_75t_R EX___U1519 ( .A(EX__n879), .Y(EX__n1191) );
  OA21x2_ASAP7_75t_R EX___U1520 ( .A1(EX__n482), .A2(EX__n990), .B(EX__n1193), .Y(EX__n1639) );
  INVx2_ASAP7_75t_R EX___U1521 ( .A(EX__n673), .Y(EX_read_reg_data_2[3]) );
  AO22x2_ASAP7_75t_R EX___U1522 ( .A1(forwarding_EX_MEM[3]), .A2(EX__n1274), .B1(
        ID_EX_read_reg_data_2[3]), .B2(EX__n480), .Y(EX__n1563) );
  INVx1_ASAP7_75t_R EX___U1523 ( .A(EX__n674), .Y(EX__n1193) );
  OA21x2_ASAP7_75t_R EX___U1524 ( .A1(EX__n1288), .A2(EX__n13), .B(EX__n1195), .Y(EX__n1613) );
  AO22x2_ASAP7_75t_R EX___U1525 ( .A1(forwarding_EX_MEM[30]), .A2(EX__n1265), .B1(
        ID_EX_read_reg_data_2[30]), .B2(EX__n423), .Y(EX__n1474) );
  INVx1_ASAP7_75t_R EX___U1526 ( .A(EX__n828), .Y(EX__n1195) );
  OA21x2_ASAP7_75t_R EX___U1527 ( .A1(EX__n1287), .A2(EX__n883), .B(EX__n1197), .Y(EX__n1615) );
  INVx2_ASAP7_75t_R EX___U1528 ( .A(EX__n676), .Y(EX_read_reg_data_2[28]) );
  AO22x2_ASAP7_75t_R EX___U1529 ( .A1(forwarding_EX_MEM[28]), .A2(EX__n1266), .B1(
        ID_EX_read_reg_data_2[28]), .B2(EX__n1263), .Y(EX__n1480) );
  INVx1_ASAP7_75t_R EX___U1530 ( .A(EX__n677), .Y(EX__n1197) );
  OA21x2_ASAP7_75t_R EX___U1531 ( .A1(EX__n1285), .A2(EX__n1134), .B(EX__n1199), .Y(EX__n1624) );
  AO22x2_ASAP7_75t_R EX___U1532 ( .A1(forwarding_EX_MEM[19]), .A2(EX__n1269), .B1(
        ID_EX_read_reg_data_2[19]), .B2(EX__n1255), .Y(EX__n1513) );
  INVx1_ASAP7_75t_R EX___U1533 ( .A(EX__n987), .Y(EX__n1199) );
  OA21x2_ASAP7_75t_R EX___U1534 ( .A1(EX__n1282), .A2(EX__n997), .B(EX__n1201), .Y(EX__n1629) );
  AO22x2_ASAP7_75t_R EX___U1535 ( .A1(forwarding_EX_MEM[14]), .A2(EX__n1270), .B1(
        ID_EX_read_reg_data_2[14]), .B2(EX__n481), .Y(EX__n1528) );
  INVx1_ASAP7_75t_R EX___U1536 ( .A(EX__n840), .Y(EX__n1201) );
  AO22x2_ASAP7_75t_R EX___U1537 ( .A1(forwarding_EX_MEM[11]), .A2(EX__n1271), .B1(
        ID_EX_read_reg_data_2[11]), .B2(EX__n1262), .Y(EX__n1536) );
  AO22x2_ASAP7_75t_R EX___U1538 ( .A1(forwarding_EX_MEM[1]), .A2(EX__n1275), .B1(
        ID_EX_read_reg_data_2[1]), .B2(EX__n1257), .Y(EX__n1568) );
  BUFx2_ASAP7_75t_R EX___U1539 ( .A(ID_EX_Branch), .Y(EX__n1204) );
  BUFx6f_ASAP7_75t_R EX___U1540 ( .A(EX__n1206), .Y(EX__n1343) );
  BUFx4f_ASAP7_75t_R EX___U1541 ( .A(EX__n1207), .Y(EX__n1206) );
  BUFx3_ASAP7_75t_R EX___U1542 ( .A(EX__n89), .Y(EX__n1207) );
  BUFx12f_ASAP7_75t_R EX___U1543 ( .A(EX__n1205), .Y(EX__n1342) );
  BUFx12f_ASAP7_75t_R EX___U1544 ( .A(EX__n1342), .Y(EX__n1341) );
  OR2x6_ASAP7_75t_R EX___U1545 ( .A(EX__n1007), .B(EX__n1008), .Y(input_A[30]) );
  OR2x6_ASAP7_75t_R EX___U1546 ( .A(EX__n1066), .B(EX__n1067), .Y(input_A[20]) );
  OR2x6_ASAP7_75t_R EX___U1547 ( .A(EX__n1098), .B(EX__n1099), .Y(input_A[26]) );
  OR2x6_ASAP7_75t_R EX___U1548 ( .A(EX__n918), .B(EX__n919), .Y(input_A[28]) );
  OR2x6_ASAP7_75t_R EX___U1549 ( .A(EX__n1158), .B(EX__n1159), .Y(input_A[27]) );
  OR2x6_ASAP7_75t_R EX___U1550 ( .A(EX__n922), .B(EX__n923), .Y(input_A[15]) );
  OR2x6_ASAP7_75t_R EX___U1551 ( .A(EX__n1070), .B(EX__n1071), .Y(input_A[16]) );
  OR2x6_ASAP7_75t_R EX___U1552 ( .A(EX__n1017), .B(EX__n1018), .Y(input_A[13]) );
  OR2x6_ASAP7_75t_R EX___U1553 ( .A(EX__n966), .B(EX__n967), .Y(input_A[14]) );
  OR2x6_ASAP7_75t_R EX___U1554 ( .A(EX__n1149), .B(EX__n1150), .Y(input_A[11]) );
  OR2x6_ASAP7_75t_R EX___U1555 ( .A(EX__n1107), .B(EX__n1108), .Y(input_A[12]) );
  OR2x6_ASAP7_75t_R EX___U1556 ( .A(EX__n927), .B(EX__n928), .Y(input_A[8]) );
  OR2x6_ASAP7_75t_R EX___U1557 ( .A(EX__n1026), .B(EX__n1027), .Y(input_A[9]) );
  OR2x6_ASAP7_75t_R EX___U1558 ( .A(EX__n971), .B(EX__n972), .Y(input_A[6]) );
  OR2x6_ASAP7_75t_R EX___U1559 ( .A(EX__n1111), .B(EX__n1112), .Y(input_A[7]) );
  OR2x6_ASAP7_75t_R EX___U1560 ( .A(EX__n1093), .B(EX__n1094), .Y(input_A[2]) );
  OR2x6_ASAP7_75t_R EX___U1561 ( .A(EX__n1058), .B(EX__n1059), .Y(input_A[3]) );
  OR2x6_ASAP7_75t_R EX___U1562 ( .A(EX__n1012), .B(EX__n1013), .Y(input_A[1]) );
  OR2x6_ASAP7_75t_R EX___U1563 ( .A(EX__n961), .B(EX__n962), .Y(input_A[0]) );
  OA22x2_ASAP7_75t_R EX___U1564 ( .A1(EX__n1210), .A2(EX__n1314), .B1(EX__n75), .B2(EX__n1209), .Y(
        input_data_2[9]) );
  INVx1_ASAP7_75t_R EX___U1565 ( .A(EX__n1544), .Y(EX__n1209) );
  INVx1_ASAP7_75t_R EX___U1566 ( .A(EX__n1545), .Y(EX__n1210) );
  OA22x2_ASAP7_75t_R EX___U1567 ( .A1(EX__n956), .A2(EX__n1310), .B1(EX__n1296), .B2(EX__n1212), 
        .Y(input_data_2[24]) );
  INVx1_ASAP7_75t_R EX___U1568 ( .A(EX__n1496), .Y(EX__n1212) );
  CKINVDCx20_ASAP7_75t_R EX___U1569 ( .A(EX__n1216), .Y(EX__n1214) );
  CKINVDCx20_ASAP7_75t_R EX___U1570 ( .A(EX__n431), .Y(EX__n1215) );
  BUFx16f_ASAP7_75t_R EX___U1571 ( .A(EX__n429), .Y(EX__n1216) );
  OR2x2_ASAP7_75t_R EX___U1572 ( .A(EX__n1325), .B(EX__n1377), .Y(EX__n1379) );
  INVx1_ASAP7_75t_R EX___U1573 ( .A(EX__n432), .Y(EX__n1217) );
  OA22x2_ASAP7_75t_R EX___U1574 ( .A1(EX__n82), .A2(EX__n989), .B1(EX__n1582), .B2(EX__n262), .Y(
        n1378) );
  INVx1_ASAP7_75t_R EX___U1575 ( .A(EX__n433), .Y(EX__n1218) );
  OR2x4_ASAP7_75t_R EX___U1576 ( .A(EX__n1217), .B(EX__n1218), .Y(input_A[29]) );
  OA22x2_ASAP7_75t_R EX___U1577 ( .A1(EX__n859), .A2(EX__n1312), .B1(EX__n70), .B2(EX__n1220), .Y(
        input_data_2[18]) );
  INVx1_ASAP7_75t_R EX___U1578 ( .A(EX__n1516), .Y(EX__n1220) );
  OA22x2_ASAP7_75t_R EX___U1579 ( .A1(EX__n812), .A2(EX__n1310), .B1(EX__n71), .B2(EX__n811), .Y(
        input_data_2[15]) );
  INVx1_ASAP7_75t_R EX___U1580 ( .A(EX__n1526), .Y(EX__n1223) );
  CKINVDCx20_ASAP7_75t_R EX___U1581 ( .A(EX__n333), .Y(EX__n1225) );
  OR2x2_ASAP7_75t_R EX___U1582 ( .A(EX__n1326), .B(EX__n1401), .Y(EX__n1403) );
  INVx1_ASAP7_75t_R EX___U1583 ( .A(EX__n334), .Y(EX__n1227) );
  OA22x2_ASAP7_75t_R EX___U1584 ( .A1(EX__n1359), .A2(EX__n752), .B1(EX__n1590), .B2(EX__n1346), 
        .Y(EX__n1402) );
  INVx1_ASAP7_75t_R EX___U1585 ( .A(EX__n335), .Y(EX__n1228) );
  OR2x4_ASAP7_75t_R EX___U1586 ( .A(EX__n1227), .B(EX__n1228), .Y(input_A[21]) );
  CKINVDCx20_ASAP7_75t_R EX___U1587 ( .A(EX__n348), .Y(EX__n1229) );
  BUFx16f_ASAP7_75t_R EX___U1588 ( .A(EX__n383), .Y(EX__n1230) );
  OR2x2_ASAP7_75t_R EX___U1589 ( .A(EX__n1331), .B(EX__n1434), .Y(EX__n1436) );
  INVx1_ASAP7_75t_R EX___U1590 ( .A(EX__n385), .Y(EX__n1231) );
  OA22x2_ASAP7_75t_R EX___U1591 ( .A1(EX__n1363), .A2(EX__n529), .B1(EX__n1601), .B2(EX__n254), .Y(
        n1435) );
  INVx1_ASAP7_75t_R EX___U1592 ( .A(EX__n386), .Y(EX__n1232) );
  OR2x4_ASAP7_75t_R EX___U1593 ( .A(EX__n1231), .B(EX__n1232), .Y(input_A[10]) );
  CKINVDCx20_ASAP7_75t_R EX___U1594 ( .A(EX__n321), .Y(EX__n1233) );
  BUFx16f_ASAP7_75t_R EX___U1595 ( .A(EX__n397), .Y(EX__n1234) );
  OR2x2_ASAP7_75t_R EX___U1596 ( .A(EX__n1334), .B(EX__n1449), .Y(EX__n1451) );
  INVx1_ASAP7_75t_R EX___U1597 ( .A(EX__n399), .Y(EX__n1235) );
  OA22x2_ASAP7_75t_R EX___U1598 ( .A1(EX__n1364), .A2(EX__n554), .B1(EX__n1080), .B2(EX__n514), .Y(
        n1450) );
  INVx1_ASAP7_75t_R EX___U1599 ( .A(EX__n400), .Y(EX__n1236) );
  OR2x4_ASAP7_75t_R EX___U1600 ( .A(EX__n1235), .B(EX__n1236), .Y(input_A[5]) );
  OR2x2_ASAP7_75t_R EX___U1601 ( .A(EX__n1324), .B(EX__n1389), .Y(EX__n1391) );
  INVx1_ASAP7_75t_R EX___U1602 ( .A(EX__n635), .Y(EX__n1240) );
  OA22x2_ASAP7_75t_R EX___U1603 ( .A1(EX__n1358), .A2(EX__n734), .B1(EX__n1081), .B2(EX__n1345), 
        .Y(EX__n1390) );
  INVx1_ASAP7_75t_R EX___U1604 ( .A(EX__n636), .Y(EX__n1241) );
  OR2x4_ASAP7_75t_R EX___U1605 ( .A(EX__n1240), .B(EX__n1241), .Y(input_A[25]) );
  OR2x2_ASAP7_75t_R EX___U1606 ( .A(EX__n1328), .B(EX__n1413), .Y(EX__n1415) );
  INVx1_ASAP7_75t_R EX___U1607 ( .A(EX__n667), .Y(EX__n1245) );
  OA22x2_ASAP7_75t_R EX___U1608 ( .A1(EX__n1360), .A2(EX__n603), .B1(EX__n1594), .B2(EX__n1347), 
        .Y(EX__n1414) );
  INVx1_ASAP7_75t_R EX___U1609 ( .A(EX__n668), .Y(EX__n1246) );
  OR2x4_ASAP7_75t_R EX___U1610 ( .A(EX__n1245), .B(EX__n1246), .Y(input_A[17]) );
  OA22x2_ASAP7_75t_R EX___U1611 ( .A1(EX__n890), .A2(EX__n1309), .B1(EX__n1306), .B2(EX__n1247), 
        .Y(input_data_2[31]) );
  INVx1_ASAP7_75t_R EX___U1612 ( .A(EX__n1472), .Y(EX__n1247) );
  INVx1_ASAP7_75t_R EX___U1613 ( .A(EX__n1473), .Y(EX__n1248) );
  BUFx12f_ASAP7_75t_R EX___U1614 ( .A(input_data_2[4]), .Y(EX__n1250) );
  OA22x2_ASAP7_75t_R EX___U1615 ( .A1(EX__n818), .A2(EX__n1315), .B1(EX__n1303), .B2(EX__n817), .Y(
        input_data_2[2]) );
  INVx1_ASAP7_75t_R EX___U1616 ( .A(EX__n1566), .Y(EX__n1253) );
  BUFx12f_ASAP7_75t_R EX___U1618 ( .A(EX__n270), .Y(EX__n1255) );
  BUFx12f_ASAP7_75t_R EX___U1619 ( .A(EX__n1259), .Y(EX__n1256) );
  BUFx12f_ASAP7_75t_R EX___U1620 ( .A(EX__n481), .Y(EX__n1257) );
  BUFx12f_ASAP7_75t_R EX___U1621 ( .A(EX__n605), .Y(EX__n1265) );
  BUFx12f_ASAP7_75t_R EX___U1622 ( .A(EX__n606), .Y(EX__n1266) );
  BUFx12f_ASAP7_75t_R EX___U1623 ( .A(EX__n1276), .Y(EX__n1275) );
  BUFx12f_ASAP7_75t_R EX___U1624 ( .A(EX__n1289), .Y(EX__n1288) );
  BUFx12f_ASAP7_75t_R EX___U1625 ( .A(EX__n308), .Y(EX__n1298) );
  BUFx12f_ASAP7_75t_R EX___U1626 ( .A(EX__n309), .Y(EX__n1299) );
  BUFx12f_ASAP7_75t_R EX___U1627 ( .A(EX__n1579), .Y(EX__n1301) );
  BUFx12f_ASAP7_75t_R EX___U1628 ( .A(EX__n1298), .Y(EX__n1302) );
  BUFx12f_ASAP7_75t_R EX___U1629 ( .A(EX__n72), .Y(EX__n1303) );
  BUFx12f_ASAP7_75t_R EX___U1630 ( .A(EX__n119), .Y(EX__n1309) );
  BUFx12f_ASAP7_75t_R EX___U1631 ( .A(EX__n120), .Y(EX__n1310) );
  BUFx12f_ASAP7_75t_R EX___U1632 ( .A(EX__n1319), .Y(EX__n1311) );
  BUFx12f_ASAP7_75t_R EX___U1633 ( .A(EX__n406), .Y(EX__n1312) );
  BUFx12f_ASAP7_75t_R EX___U1634 ( .A(EX__n407), .Y(EX__n1313) );
  BUFx12f_ASAP7_75t_R EX___U1635 ( .A(EX__n458), .Y(EX__n1344) );
  BUFx12f_ASAP7_75t_R EX___U1636 ( .A(EX__n1350), .Y(EX__n1348) );
  BUFx12f_ASAP7_75t_R EX___U1637 ( .A(EX__n1355), .Y(EX__n1349) );
  BUFx12f_ASAP7_75t_R EX___U1638 ( .A(EX__n1351), .Y(EX__n1350) );
  BUFx12f_ASAP7_75t_R EX___U1639 ( .A(EX__n517), .Y(EX__n1356) );
  BUFx12f_ASAP7_75t_R EX___U1640 ( .A(EX__n518), .Y(EX__n1357) );
  BUFx12f_ASAP7_75t_R EX___U1641 ( .A(EX__n101), .Y(EX__n1365) );
  INVx1_ASAP7_75t_R EX___U1642 ( .A(forwarding_EX_MEM[31]), .Y(EX__n1371) );
  INVx1_ASAP7_75t_R EX___U1643 ( .A(forwarding_EX_MEM[30]), .Y(EX__n1374) );
  INVx1_ASAP7_75t_R EX___U1644 ( .A(forwarding_EX_MEM[29]), .Y(EX__n1377) );
  INVx1_ASAP7_75t_R EX___U1645 ( .A(forwarding_EX_MEM[28]), .Y(EX__n1380) );
  INVx1_ASAP7_75t_R EX___U1646 ( .A(forwarding_EX_MEM[27]), .Y(EX__n1383) );
  INVx1_ASAP7_75t_R EX___U1647 ( .A(forwarding_EX_MEM[26]), .Y(EX__n1386) );
  INVx1_ASAP7_75t_R EX___U1648 ( .A(forwarding_EX_MEM[25]), .Y(EX__n1389) );
  INVx1_ASAP7_75t_R EX___U1649 ( .A(forwarding_EX_MEM[24]), .Y(EX__n1392) );
  INVx1_ASAP7_75t_R EX___U1650 ( .A(forwarding_EX_MEM[23]), .Y(EX__n1395) );
  INVx1_ASAP7_75t_R EX___U1651 ( .A(forwarding_EX_MEM[22]), .Y(EX__n1398) );
  INVx1_ASAP7_75t_R EX___U1652 ( .A(forwarding_EX_MEM[21]), .Y(EX__n1401) );
  INVx1_ASAP7_75t_R EX___U1653 ( .A(forwarding_EX_MEM[20]), .Y(EX__n1404) );
  INVx1_ASAP7_75t_R EX___U1654 ( .A(forwarding_EX_MEM[19]), .Y(EX__n1407) );
  INVx1_ASAP7_75t_R EX___U1655 ( .A(forwarding_EX_MEM[18]), .Y(EX__n1410) );
  INVx1_ASAP7_75t_R EX___U1656 ( .A(forwarding_EX_MEM[17]), .Y(EX__n1413) );
  INVx1_ASAP7_75t_R EX___U1657 ( .A(forwarding_EX_MEM[16]), .Y(EX__n1416) );
  INVx1_ASAP7_75t_R EX___U1658 ( .A(forwarding_EX_MEM[15]), .Y(EX__n1419) );
  INVx1_ASAP7_75t_R EX___U1659 ( .A(forwarding_EX_MEM[14]), .Y(EX__n1422) );
  INVx1_ASAP7_75t_R EX___U1660 ( .A(forwarding_EX_MEM[13]), .Y(EX__n1425) );
  INVx1_ASAP7_75t_R EX___U1661 ( .A(forwarding_EX_MEM[12]), .Y(EX__n1428) );
  INVx1_ASAP7_75t_R EX___U1662 ( .A(forwarding_EX_MEM[11]), .Y(EX__n1431) );
  INVx1_ASAP7_75t_R EX___U1663 ( .A(forwarding_EX_MEM[10]), .Y(EX__n1434) );
  INVx1_ASAP7_75t_R EX___U1664 ( .A(forwarding_EX_MEM[9]), .Y(EX__n1437) );
  INVx1_ASAP7_75t_R EX___U1665 ( .A(forwarding_EX_MEM[8]), .Y(EX__n1440) );
  INVx1_ASAP7_75t_R EX___U1666 ( .A(forwarding_EX_MEM[7]), .Y(EX__n1443) );
  INVx1_ASAP7_75t_R EX___U1667 ( .A(forwarding_EX_MEM[6]), .Y(EX__n1446) );
  INVx1_ASAP7_75t_R EX___U1668 ( .A(forwarding_EX_MEM[5]), .Y(EX__n1449) );
  INVx1_ASAP7_75t_R EX___U1669 ( .A(forwarding_EX_MEM[4]), .Y(EX__n1452) );
  INVx1_ASAP7_75t_R EX___U1670 ( .A(forwarding_EX_MEM[3]), .Y(EX__n1455) );
  INVx1_ASAP7_75t_R EX___U1671 ( .A(forwarding_EX_MEM[2]), .Y(EX__n1458) );
  INVx1_ASAP7_75t_R EX___U1672 ( .A(forwarding_EX_MEM[1]), .Y(EX__n1461) );
  INVx1_ASAP7_75t_R EX___U1673 ( .A(forwarding_EX_MEM[0]), .Y(EX__n1464) );
  INVx1_ASAP7_75t_R EX___U1674 ( .A(ForwardB[1]), .Y(EX__n1467) );
  INVx1_ASAP7_75t_R EX___U1675 ( .A(ForwardB[0]), .Y(EX__n1468) );
  INVx1_ASAP7_75t_R EX___U1676 ( .A(ID_EX_imm[23]), .Y(EX__n1499) );
  INVx1_ASAP7_75t_R EX___U1677 ( .A(ID_EX_imm[21]), .Y(EX__n1507) );
  AND2x2_ASAP7_75t_R EX___U1678 ( .A(EX__n1204), .B(EX__n1148), .Y(EX__n1641) );
  INVx1_ASAP7_75t_R EX___U1679 ( .A(ID_EX_read_reg_data_1[31]), .Y(EX__n1580) );
  INVx1_ASAP7_75t_R EX___U1680 ( .A(ID_EX_read_reg_data_1[30]), .Y(EX__n1581) );
  INVx1_ASAP7_75t_R EX___U1681 ( .A(ID_EX_read_reg_data_1[29]), .Y(EX__n1582) );
  INVx1_ASAP7_75t_R EX___U1682 ( .A(ID_EX_read_reg_data_1[28]), .Y(EX__n1583) );
  INVx1_ASAP7_75t_R EX___U1683 ( .A(ID_EX_read_reg_data_1[27]), .Y(EX__n1584) );
  INVx1_ASAP7_75t_R EX___U1684 ( .A(ID_EX_read_reg_data_1[26]), .Y(EX__n1585) );
  INVx1_ASAP7_75t_R EX___U1685 ( .A(ID_EX_read_reg_data_1[24]), .Y(EX__n1587) );
  INVx1_ASAP7_75t_R EX___U1686 ( .A(ID_EX_read_reg_data_1[21]), .Y(EX__n1590) );
  INVx1_ASAP7_75t_R EX___U1687 ( .A(ID_EX_read_reg_data_1[20]), .Y(EX__n1591) );
  INVx1_ASAP7_75t_R EX___U1688 ( .A(ID_EX_read_reg_data_1[19]), .Y(EX__n1592) );
  INVx1_ASAP7_75t_R EX___U1689 ( .A(ID_EX_read_reg_data_1[18]), .Y(EX__n1593) );
  INVx1_ASAP7_75t_R EX___U1690 ( .A(ID_EX_read_reg_data_1[17]), .Y(EX__n1594) );
  INVx1_ASAP7_75t_R EX___U1691 ( .A(ID_EX_read_reg_data_1[16]), .Y(EX__n1595) );
  INVx1_ASAP7_75t_R EX___U1692 ( .A(ID_EX_read_reg_data_1[15]), .Y(EX__n1596) );
  INVx1_ASAP7_75t_R EX___U1693 ( .A(ID_EX_read_reg_data_1[14]), .Y(EX__n1597) );
  INVx1_ASAP7_75t_R EX___U1694 ( .A(ID_EX_read_reg_data_1[13]), .Y(EX__n1598) );
  INVx1_ASAP7_75t_R EX___U1695 ( .A(ID_EX_read_reg_data_1[12]), .Y(EX__n1599) );
  INVx1_ASAP7_75t_R EX___U1696 ( .A(ID_EX_read_reg_data_1[10]), .Y(EX__n1601) );
  INVx1_ASAP7_75t_R EX___U1697 ( .A(ID_EX_read_reg_data_1[9]), .Y(EX__n1602) );
  INVx1_ASAP7_75t_R EX___U1698 ( .A(ID_EX_read_reg_data_1[8]), .Y(EX__n1603) );
  INVx1_ASAP7_75t_R EX___U1699 ( .A(ID_EX_read_reg_data_1[7]), .Y(EX__n1604) );
  INVx1_ASAP7_75t_R EX___U1700 ( .A(ID_EX_read_reg_data_1[6]), .Y(EX__n1605) );
  INVx1_ASAP7_75t_R EX___U1701 ( .A(ID_EX_read_reg_data_1[4]), .Y(EX__n1607) );
  INVx1_ASAP7_75t_R EX___U1702 ( .A(ID_EX_read_reg_data_1[3]), .Y(EX__n1608) );
  INVx1_ASAP7_75t_R EX___U1703 ( .A(ID_EX_read_reg_data_1[2]), .Y(EX__n1609) );
  INVx1_ASAP7_75t_R EX___U1704 ( .A(ID_EX_read_reg_data_1[1]), .Y(EX__n1610) );
  INVx1_ASAP7_75t_R EX___U1705 ( .A(ID_EX_read_reg_data_1[0]), .Y(EX__n1611) );
  
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___MemWrite_out_reg ( .D(EX_MEM__n280), .CLK(clk), .SETN(EX_MEM__EX_MEM__n145), 
        .RESETN(EX_MEM__n14), .QN(EX_MEM_MemWrite) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___rd_out_reg_4_ ( .D(EX_MEM__n273), .CLK(clk), .SETN(EX_MEM__EX_MEM__n145), 
        .RESETN(EX_MEM__n14), .QN(EX_MEM__n316) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___rd_out_reg_3_ ( .D(EX_MEM__n274), .CLK(clk), .SETN(EX_MEM__EX_MEM__n145), 
        .RESETN(EX_MEM__n14), .QN(EX_MEM__n317) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___rd_out_reg_2_ ( .D(EX_MEM__n275), .CLK(clk), .SETN(EX_MEM__EX_MEM__n145), 
        .RESETN(EX_MEM__n14), .QN(EX_MEM__n318) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___rd_out_reg_1_ ( .D(EX_MEM__n276), .CLK(clk), .SETN(EX_MEM__EX_MEM__n145), 
        .RESETN(EX_MEM__n14), .QN(EX_MEM__n319) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___rd_out_reg_0_ ( .D(EX_MEM__n277), .CLK(clk), .SETN(EX_MEM__EX_MEM__n145), 
        .RESETN(EX_MEM__n14), .QN(EX_MEM__n320) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___RegWrite_out_reg ( .D(EX_MEM__n127), .CLK(clk), .SETN(EX_MEM__EX_MEM__n145), 
        .RESETN(EX_MEM__n14), .QN(EX_MEM__n283) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_31_ ( .D(EX_MEM__n129), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n284) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_30_ ( .D(EX_MEM__n77), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n285) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_29_ ( .D(EX_MEM__n49), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n286) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_28_ ( .D(EX_MEM__n73), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n287) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_27_ ( .D(EX_MEM__n118), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n288) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_26_ ( .D(EX_MEM__n119), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n289) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_25_ ( .D(EX_MEM__n78), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n290) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_24_ ( .D(EX_MEM__n79), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n291) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_23_ ( .D(EX_MEM__n120), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n292) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_22_ ( .D(EX_MEM__n121), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n293) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_21_ ( .D(EX_MEM__n80), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n294) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_20_ ( .D(EX_MEM__n122), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n295) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_19_ ( .D(EX_MEM__n42), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n296) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_18_ ( .D(EX_MEM__n25), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n297) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_17_ ( .D(EX_MEM__n43), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n298) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_16_ ( .D(EX_MEM__n123), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n299) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_15_ ( .D(EX_MEM__n124), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n300) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_14_ ( .D(EX_MEM__n81), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n301) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_13_ ( .D(EX_MEM__n125), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n302) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_12_ ( .D(EX_MEM__n44), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n303) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_11_ ( .D(EX_MEM__n45), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n304) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_10_ ( .D(EX_MEM__n46), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n305) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_9_ ( .D(EX_MEM__n74), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n306) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_8_ ( .D(EX_MEM__n75), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n307) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_7_ ( .D(EX_MEM__n250), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n308) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_6_ ( .D(EX_MEM__n130), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n309) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_5_ ( .D(EX_MEM__n76), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n310) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_4_ ( .D(EX_MEM__n131), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n311) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_3_ ( .D(EX_MEM__n254), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n312) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_2_ ( .D(EX_MEM__n126), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n313) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_1_ ( .D(EX_MEM__n47), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n314) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___ALU_result_out_reg_0_ ( .D(EX_MEM__n48), .CLK(clk), .SETN(
        EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM__n315) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_29_ ( .D(EX_MEM__n36), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[29]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_28_ ( .D(EX_MEM__n69), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[28]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_27_ ( .D(EX_MEM__n10), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[27]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_26_ ( .D(EX_MEM__n70), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[26]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_25_ ( .D(EX_MEM__n1), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[25]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_24_ ( .D(EX_MEM__n5), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[24]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_23_ ( .D(EX_MEM__n265), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[23]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_22_ ( .D(EX_MEM__n264), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[22]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_21_ ( .D(EX_MEM__n71), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[21]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_20_ ( .D(EX_MEM__n37), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[20]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_19_ ( .D(EX_MEM__n41), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[19]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_18_ ( .D(EX_MEM__n4), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[18]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_17_ ( .D(EX_MEM__n260), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[17]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_16_ ( .D(EX_MEM__n6), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[16]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_15_ ( .D(EX_MEM__n3), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[15]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_14_ ( .D(EX_MEM__n259), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[14]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_13_ ( .D(EX_MEM__n258), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[13]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_11_ ( .D(EX_MEM__n8), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[11]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_10_ ( .D(EX_MEM__n13), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[10]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_9_ ( .D(EX_MEM__n12), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[9]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_8_ ( .D(EX_MEM__n72), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[8]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_7_ ( .D(EX_MEM__n7), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[7]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_6_ ( .D(EX_MEM__n2), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[6]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_5_ ( .D(EX_MEM__n270), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[5]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_4_ ( .D(EX_MEM__n132), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[4]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_3_ ( .D(EX_MEM__n16), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[3]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_2_ ( .D(EX_MEM__n38), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[2]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_1_ ( .D(EX_MEM__n40), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[1]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_0_ ( .D(EX_MEM__n39), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[0]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___MemRead_out_reg ( .D(EX_MEM__n35), .CLK(clk), .SETN(EX_MEM__EX_MEM__n145), 
        .RESETN(EX_MEM__n14), .QN(EX_MEM__n281) );
  CKINVDCx10_ASAP7_75t_R EX_MEM___U147 ( .A(rst), .Y(EX_MEM__n145) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___MemtoReg_out_reg ( .D(EX_MEM__n279), .CLK(clk), .SETN(EX_MEM__EX_MEM__n145), 
        .RESETN(EX_MEM__n14), .QN(EX_MEM__n282) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_12_ ( .D(EX_MEM__n15), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[12]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_31_ ( .D(EX_MEM__n268), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[31]) );
  DFFASRHQNx1_ASAP7_75t_R EX_MEM___read_reg_data_2_out_reg_30_ ( .D(EX_MEM__n267), .CLK(clk), 
        .SETN(EX_MEM__EX_MEM__n145), .RESETN(EX_MEM__n14), .QN(EX_MEM_read_reg_data_2[30]) );
  TIEHIx1_ASAP7_75t_R EX_MEM___U3 ( .H(EX_MEM__n14) );
  HB1xp67_ASAP7_75t_R EX_MEM___U4 ( .A(EX_read_reg_data_2[21]), .Y(EX_MEM__n263) );
  INVx1_ASAP7_75t_R EX_MEM___U5 ( .A(EX_MEM__n263), .Y(EX_MEM__n71) );
  INVxp67_ASAP7_75t_R EX_MEM___U6 ( .A(EX_read_reg_data_2[23]), .Y(EX_MEM__n265) );
  INVxp67_ASAP7_75t_R EX_MEM___U7 ( .A(EX_MEM__n266), .Y(EX_MEM__n70) );
  HB1xp67_ASAP7_75t_R EX_MEM___U8 ( .A(EX_read_reg_data_2[26]), .Y(EX_MEM__n266) );
  INVx1_ASAP7_75t_R EX_MEM___U9 ( .A(n18), .Y(EX_MEM__n267) );
  INVxp33_ASAP7_75t_R EX_MEM___U10 ( .A(ID_EX_rd[2]), .Y(EX_MEM__n275) );
  INVxp67_ASAP7_75t_R EX_MEM___U11 ( .A(EX_read_reg_data_2[24]), .Y(EX_MEM__n5) );
  INVx1_ASAP7_75t_R EX_MEM___U12 ( .A(EX_read_reg_data_2[25]), .Y(EX_MEM__n1) );
  INVx1_ASAP7_75t_R EX_MEM___U13 ( .A(EX_read_reg_data_2[6]), .Y(EX_MEM__n2) );
  INVxp67_ASAP7_75t_R EX_MEM___U14 ( .A(n20), .Y(EX_MEM__n3) );
  HB1xp67_ASAP7_75t_R EX_MEM___U15 ( .A(EX_MEM__n309), .Y(EX_MEM__n109) );
  INVxp67_ASAP7_75t_R EX_MEM___U16 ( .A(EX_read_reg_data_2[18]), .Y(EX_MEM__n4) );
  INVxp67_ASAP7_75t_R EX_MEM___U17 ( .A(EX_read_reg_data_2[5]), .Y(EX_MEM__n270) );
  INVxp67_ASAP7_75t_R EX_MEM___U18 ( .A(EX_read_reg_data_2[12]), .Y(EX_MEM__n15) );
  INVx1_ASAP7_75t_R EX_MEM___U19 ( .A(EX_read_reg_data_2[16]), .Y(EX_MEM__n6) );
  INVx1_ASAP7_75t_R EX_MEM___U20 ( .A(EX_read_reg_data_2[7]), .Y(EX_MEM__n7) );
  INVxp33_ASAP7_75t_R EX_MEM___U21 ( .A(EX_read_reg_data_2[29]), .Y(EX_MEM__n9) );
  INVx1_ASAP7_75t_R EX_MEM___U22 ( .A(EX_read_reg_data_2[11]), .Y(EX_MEM__n8) );
  INVx2_ASAP7_75t_R EX_MEM___U23 ( .A(EX_MEM__n271), .Y(EX_MEM__n72) );
  BUFx3_ASAP7_75t_R EX_MEM___U24 ( .A(EX_read_reg_data_2[8]), .Y(EX_MEM__n271) );
  INVx1_ASAP7_75t_R EX_MEM___U25 ( .A(EX_read_reg_data_2[27]), .Y(EX_MEM__n10) );
  INVxp33_ASAP7_75t_R EX_MEM___U26 ( .A(EX_read_reg_data_2[0]), .Y(EX_MEM__n11) );
  HB1xp67_ASAP7_75t_R EX_MEM___U27 ( .A(EX_MEM__n9), .Y(EX_MEM__n36) );
  INVxp67_ASAP7_75t_R EX_MEM___U28 ( .A(EX_MEM__n269), .Y(EX_MEM__n16) );
  HB1xp67_ASAP7_75t_R EX_MEM___U29 ( .A(EX_read_reg_data_2[3]), .Y(EX_MEM__n269) );
  INVxp67_ASAP7_75t_R EX_MEM___U30 ( .A(EX_read_reg_data_2[28]), .Y(EX_MEM__n69) );
  HB1xp67_ASAP7_75t_R EX_MEM___U31 ( .A(EX_MEM__n133), .Y(EX_MEM__n38) );
  INVxp33_ASAP7_75t_R EX_MEM___U32 ( .A(EX_read_reg_data_2[2]), .Y(EX_MEM__n133) );
  INVx1_ASAP7_75t_R EX_MEM___U33 ( .A(EX_read_reg_data_2[9]), .Y(EX_MEM__n12) );
  INVxp67_ASAP7_75t_R EX_MEM___U34 ( .A(EX_MEM__n261), .Y(EX_MEM__n40) );
  HB1xp67_ASAP7_75t_R EX_MEM___U35 ( .A(EX_read_reg_data_2[1]), .Y(EX_MEM__n261) );
  INVxp67_ASAP7_75t_R EX_MEM___U36 ( .A(EX_read_reg_data_2[19]), .Y(EX_MEM__n41) );
  INVx1_ASAP7_75t_R EX_MEM___U37 ( .A(EX_read_reg_data_2[10]), .Y(EX_MEM__n13) );
  HB1xp67_ASAP7_75t_R EX_MEM___U38 ( .A(EX_MEM__n134), .Y(EX_MEM__n37) );
  INVxp33_ASAP7_75t_R EX_MEM___U39 ( .A(EX_MEM__n262), .Y(EX_MEM__n134) );
  HB1xp67_ASAP7_75t_R EX_MEM___U40 ( .A(EX_MEM__n11), .Y(EX_MEM__n39) );
  HB1xp67_ASAP7_75t_R EX_MEM___U41 ( .A(EX_read_reg_data_2[20]), .Y(EX_MEM__n262) );
  BUFx6f_ASAP7_75t_R EX_MEM___U42 ( .A(EX_MEM__n117), .Y(EX_MEM_RegWrite) );
  BUFx3_ASAP7_75t_R EX_MEM___U43 ( .A(EX_MEM__n18), .Y(EX_MEM__n17) );
  BUFx2_ASAP7_75t_R EX_MEM___U44 ( .A(EX_MEM__n317), .Y(EX_MEM__n18) );
  BUFx12f_ASAP7_75t_R EX_MEM___U45 ( .A(EX_MEM__n20), .Y(EX_MEM__n19) );
  BUFx12f_ASAP7_75t_R EX_MEM___U46 ( .A(EX_MEM__n219), .Y(EX_MEM__n20) );
  BUFx3_ASAP7_75t_R EX_MEM___U47 ( .A(EX_MEM__n22), .Y(EX_MEM__n21) );
  BUFx2_ASAP7_75t_R EX_MEM___U48 ( .A(EX_MEM__n320), .Y(EX_MEM__n22) );
  BUFx12f_ASAP7_75t_R EX_MEM___U49 ( .A(EX_MEM__n24), .Y(EX_MEM__n23) );
  BUFx12f_ASAP7_75t_R EX_MEM___U50 ( .A(EX_MEM__n225), .Y(EX_MEM__n24) );
  BUFx2_ASAP7_75t_R EX_MEM___U51 ( .A(EX_ALU_result[18]), .Y(EX_MEM__n239) );
  INVx1_ASAP7_75t_R EX_MEM___U52 ( .A(EX_MEM__n239), .Y(EX_MEM__n25) );
  BUFx3_ASAP7_75t_R EX_MEM___U53 ( .A(EX_MEM__n27), .Y(EX_MEM__n26) );
  BUFx2_ASAP7_75t_R EX_MEM___U54 ( .A(EX_MEM__n316), .Y(EX_MEM__n27) );
  BUFx12f_ASAP7_75t_R EX_MEM___U55 ( .A(EX_MEM__n29), .Y(EX_MEM__n28) );
  BUFx12f_ASAP7_75t_R EX_MEM___U56 ( .A(EX_MEM__n217), .Y(EX_MEM__n29) );
  BUFx3_ASAP7_75t_R EX_MEM___U57 ( .A(EX_MEM__n31), .Y(EX_MEM__n30) );
  BUFx2_ASAP7_75t_R EX_MEM___U58 ( .A(EX_MEM__EX_MEM__n318), .Y(EX_MEM__n31) );
  BUFx12f_ASAP7_75t_R EX_MEM___U59 ( .A(EX_MEM__n33), .Y(EX_MEM__n32) );
  BUFx12f_ASAP7_75t_R EX_MEM___U60 ( .A(EX_MEM__n221), .Y(EX_MEM__n33) );
  BUFx12f_ASAP7_75t_R EX_MEM___U61 ( .A(EX_MEM__n319), .Y(EX_MEM__n34) );
  BUFx2_ASAP7_75t_R EX_MEM___U62 ( .A(EX_MEM__n128), .Y(EX_MEM__n35) );
  BUFx2_ASAP7_75t_R EX_MEM___U63 ( .A(EX_ALU_result[19]), .Y(EX_MEM__n238) );
  INVx1_ASAP7_75t_R EX_MEM___U64 ( .A(EX_MEM__n238), .Y(EX_MEM__n42) );
  BUFx2_ASAP7_75t_R EX_MEM___U65 ( .A(EX_ALU_result[17]), .Y(EX_MEM__n240) );
  INVx1_ASAP7_75t_R EX_MEM___U66 ( .A(EX_MEM__n240), .Y(EX_MEM__n43) );
  BUFx2_ASAP7_75t_R EX_MEM___U67 ( .A(EX_ALU_result[12]), .Y(EX_MEM__n245) );
  INVx1_ASAP7_75t_R EX_MEM___U68 ( .A(EX_MEM__n245), .Y(EX_MEM__n44) );
  BUFx2_ASAP7_75t_R EX_MEM___U69 ( .A(EX_ALU_result[11]), .Y(EX_MEM__n246) );
  INVx1_ASAP7_75t_R EX_MEM___U70 ( .A(EX_MEM__n246), .Y(EX_MEM__n45) );
  BUFx2_ASAP7_75t_R EX_MEM___U71 ( .A(EX_ALU_result[10]), .Y(EX_MEM__n247) );
  INVx1_ASAP7_75t_R EX_MEM___U72 ( .A(EX_MEM__n247), .Y(EX_MEM__n46) );
  BUFx2_ASAP7_75t_R EX_MEM___U73 ( .A(EX_ALU_result[1]), .Y(EX_MEM__n256) );
  INVx1_ASAP7_75t_R EX_MEM___U74 ( .A(EX_MEM__n256), .Y(EX_MEM__n47) );
  BUFx2_ASAP7_75t_R EX_MEM___U75 ( .A(EX_ALU_result[0]), .Y(EX_MEM__n257) );
  INVx1_ASAP7_75t_R EX_MEM___U76 ( .A(EX_MEM__n257), .Y(EX_MEM__n48) );
  BUFx2_ASAP7_75t_R EX_MEM___U77 ( .A(EX_ALU_result[29]), .Y(EX_MEM__n228) );
  INVx1_ASAP7_75t_R EX_MEM___U78 ( .A(EX_MEM__n228), .Y(EX_MEM__n49) );
  BUFx2_ASAP7_75t_R EX_MEM___U79 ( .A(EX_MEM__n283), .Y(EX_MEM__n50) );
  BUFx3_ASAP7_75t_R EX_MEM___U80 ( .A(EX_MEM__n52), .Y(EX_MEM__n51) );
  BUFx2_ASAP7_75t_R EX_MEM___U81 ( .A(EX_MEM__n284), .Y(EX_MEM__n52) );
  BUFx3_ASAP7_75t_R EX_MEM___U82 ( .A(EX_MEM__n54), .Y(EX_MEM__n53) );
  BUFx2_ASAP7_75t_R EX_MEM___U83 ( .A(EX_MEM__n289), .Y(EX_MEM__n54) );
  BUFx3_ASAP7_75t_R EX_MEM___U84 ( .A(EX_MEM__n56), .Y(EX_MEM__n55) );
  BUFx2_ASAP7_75t_R EX_MEM___U85 ( .A(EX_MEM__n290), .Y(EX_MEM__n56) );
  BUFx3_ASAP7_75t_R EX_MEM___U86 ( .A(EX_MEM__n58), .Y(EX_MEM__n57) );
  BUFx2_ASAP7_75t_R EX_MEM___U87 ( .A(EX_MEM__n294), .Y(EX_MEM__n58) );
  BUFx3_ASAP7_75t_R EX_MEM___U88 ( .A(EX_MEM__n60), .Y(EX_MEM__n59) );
  BUFx2_ASAP7_75t_R EX_MEM___U89 ( .A(EX_MEM__n297), .Y(EX_MEM__n60) );
  BUFx3_ASAP7_75t_R EX_MEM___U90 ( .A(EX_MEM__n62), .Y(EX_MEM__n61) );
  BUFx2_ASAP7_75t_R EX_MEM___U91 ( .A(EX_MEM__n308), .Y(EX_MEM__n62) );
  BUFx3_ASAP7_75t_R EX_MEM___U92 ( .A(EX_MEM__n64), .Y(EX_MEM__n63) );
  BUFx2_ASAP7_75t_R EX_MEM___U93 ( .A(EX_MEM__n310), .Y(EX_MEM__n64) );
  BUFx3_ASAP7_75t_R EX_MEM___U94 ( .A(EX_MEM__n66), .Y(EX_MEM__n65) );
  BUFx2_ASAP7_75t_R EX_MEM___U95 ( .A(EX_MEM__n311), .Y(EX_MEM__n66) );
  BUFx3_ASAP7_75t_R EX_MEM___U96 ( .A(EX_MEM__n68), .Y(EX_MEM__n67) );
  BUFx2_ASAP7_75t_R EX_MEM___U97 ( .A(EX_MEM__n313), .Y(EX_MEM__n68) );
  BUFx12f_ASAP7_75t_R EX_MEM___U98 ( .A(EX_MEM__n23), .Y(EX_MEM_rd[0]) );
  BUFx2_ASAP7_75t_R EX_MEM___U99 ( .A(EX_ALU_result[28]), .Y(EX_MEM__n229) );
  INVx1_ASAP7_75t_R EX_MEM___U100 ( .A(EX_MEM__n229), .Y(EX_MEM__n73) );
  BUFx2_ASAP7_75t_R EX_MEM___U101 ( .A(EX_ALU_result[9]), .Y(EX_MEM__n248) );
  INVx1_ASAP7_75t_R EX_MEM___U102 ( .A(EX_MEM__n248), .Y(EX_MEM__n74) );
  BUFx2_ASAP7_75t_R EX_MEM___U103 ( .A(EX_ALU_result[8]), .Y(EX_MEM__n249) );
  INVx1_ASAP7_75t_R EX_MEM___U104 ( .A(EX_MEM__n249), .Y(EX_MEM__n75) );
  BUFx2_ASAP7_75t_R EX_MEM___U105 ( .A(EX_ALU_result[5]), .Y(EX_MEM__n252) );
  INVx1_ASAP7_75t_R EX_MEM___U106 ( .A(EX_MEM__n252), .Y(EX_MEM__n76) );
  BUFx2_ASAP7_75t_R EX_MEM___U107 ( .A(EX_ALU_result[30]), .Y(EX_MEM__n227) );
  INVx1_ASAP7_75t_R EX_MEM___U108 ( .A(EX_MEM__n227), .Y(EX_MEM__n77) );
  BUFx2_ASAP7_75t_R EX_MEM___U109 ( .A(EX_MEM__n232), .Y(EX_MEM__n78) );
  BUFx2_ASAP7_75t_R EX_MEM___U110 ( .A(EX_MEM__n233), .Y(EX_MEM__n79) );
  BUFx2_ASAP7_75t_R EX_MEM___U111 ( .A(EX_ALU_result[21]), .Y(EX_MEM__n236) );
  INVx1_ASAP7_75t_R EX_MEM___U112 ( .A(EX_MEM__n236), .Y(EX_MEM__n80) );
  BUFx2_ASAP7_75t_R EX_MEM___U113 ( .A(EX_ALU_result[14]), .Y(EX_MEM__n243) );
  INVx1_ASAP7_75t_R EX_MEM___U114 ( .A(EX_MEM__n243), .Y(EX_MEM__n81) );
  BUFx2_ASAP7_75t_R EX_MEM___U115 ( .A(EX_MEM__n83), .Y(EX_MEM_MemRead) );
  BUFx2_ASAP7_75t_R EX_MEM___U116 ( .A(EX_MEM__n281), .Y(EX_MEM__n83) );
  BUFx2_ASAP7_75t_R EX_MEM___U117 ( .A(EX_MEM__n85), .Y(EX_MEM_MemToReg) );
  BUFx2_ASAP7_75t_R EX_MEM___U118 ( .A(EX_MEM__n282), .Y(EX_MEM__n85) );
  BUFx3_ASAP7_75t_R EX_MEM___U119 ( .A(EX_MEM__n87), .Y(EX_MEM__n86) );
  BUFx2_ASAP7_75t_R EX_MEM___U120 ( .A(EX_MEM__n286), .Y(EX_MEM__n87) );
  BUFx3_ASAP7_75t_R EX_MEM___U121 ( .A(EX_MEM__n89), .Y(EX_MEM__n88) );
  BUFx2_ASAP7_75t_R EX_MEM___U122 ( .A(EX_MEM__n288), .Y(EX_MEM__n89) );
  BUFx3_ASAP7_75t_R EX_MEM___U123 ( .A(EX_MEM__n91), .Y(EX_MEM__n90) );
  BUFx2_ASAP7_75t_R EX_MEM___U124 ( .A(EX_MEM__n292), .Y(EX_MEM__n91) );
  BUFx3_ASAP7_75t_R EX_MEM___U125 ( .A(EX_MEM__n93), .Y(EX_MEM__n92) );
  BUFx2_ASAP7_75t_R EX_MEM___U126 ( .A(EX_MEM__n293), .Y(EX_MEM__n93) );
  BUFx3_ASAP7_75t_R EX_MEM___U127 ( .A(EX_MEM__n95), .Y(EX_MEM__n94) );
  BUFx2_ASAP7_75t_R EX_MEM___U128 ( .A(EX_MEM__n295), .Y(EX_MEM__n95) );
  BUFx3_ASAP7_75t_R EX_MEM___U129 ( .A(EX_MEM__n97), .Y(EX_MEM__n96) );
  BUFx2_ASAP7_75t_R EX_MEM___U130 ( .A(EX_MEM__n298), .Y(EX_MEM__n97) );
  BUFx3_ASAP7_75t_R EX_MEM___U131 ( .A(EX_MEM__n99), .Y(EX_MEM__n98) );
  BUFx2_ASAP7_75t_R EX_MEM___U132 ( .A(EX_MEM__n299), .Y(EX_MEM__n99) );
  BUFx3_ASAP7_75t_R EX_MEM___U133 ( .A(EX_MEM__n101), .Y(EX_MEM__n100) );
  BUFx2_ASAP7_75t_R EX_MEM___U134 ( .A(EX_MEM__n300), .Y(EX_MEM__n101) );
  BUFx3_ASAP7_75t_R EX_MEM___U135 ( .A(EX_MEM__n103), .Y(EX_MEM__n102) );
  BUFx2_ASAP7_75t_R EX_MEM___U136 ( .A(EX_MEM__n302), .Y(EX_MEM__n103) );
  BUFx3_ASAP7_75t_R EX_MEM___U137 ( .A(EX_MEM__n105), .Y(EX_MEM__n104) );
  BUFx2_ASAP7_75t_R EX_MEM___U138 ( .A(EX_MEM__n304), .Y(EX_MEM__n105) );
  BUFx3_ASAP7_75t_R EX_MEM___U139 ( .A(EX_MEM__n107), .Y(EX_MEM__n106) );
  BUFx2_ASAP7_75t_R EX_MEM___U140 ( .A(EX_MEM__n305), .Y(EX_MEM__n107) );
  BUFx3_ASAP7_75t_R EX_MEM___U141 ( .A(EX_MEM__n109), .Y(EX_MEM__n108) );
  BUFx3_ASAP7_75t_R EX_MEM___U142 ( .A(EX_MEM__n111), .Y(EX_MEM__n110) );
  BUFx2_ASAP7_75t_R EX_MEM___U143 ( .A(EX_MEM__n312), .Y(EX_MEM__n111) );
  BUFx3_ASAP7_75t_R EX_MEM___U144 ( .A(EX_MEM__n113), .Y(EX_MEM__n112) );
  BUFx2_ASAP7_75t_R EX_MEM___U145 ( .A(EX_MEM__n314), .Y(EX_MEM__n113) );
  BUFx3_ASAP7_75t_R EX_MEM___U146 ( .A(EX_MEM__n115), .Y(EX_MEM__n114) );
  BUFx2_ASAP7_75t_R EX_MEM___U148 ( .A(EX_MEM__n315), .Y(EX_MEM__n115) );
  BUFx3_ASAP7_75t_R EX_MEM___U149 ( .A(EX_MEM__n50), .Y(EX_MEM__n117) );
  BUFx12f_ASAP7_75t_R EX_MEM___U150 ( .A(EX_MEM__n19), .Y(EX_MEM_rd[3]) );
  BUFx12f_ASAP7_75t_R EX_MEM___U151 ( .A(EX_MEM__n28), .Y(EX_MEM_rd[4]) );
  BUFx2_ASAP7_75t_R EX_MEM___U152 ( .A(EX_MEM__n230), .Y(EX_MEM__n118) );
  BUFx2_ASAP7_75t_R EX_MEM___U153 ( .A(EX_MEM__n231), .Y(EX_MEM__n119) );
  BUFx2_ASAP7_75t_R EX_MEM___U154 ( .A(EX_ALU_result[23]), .Y(EX_MEM__n234) );
  INVx1_ASAP7_75t_R EX_MEM___U155 ( .A(EX_MEM__n234), .Y(EX_MEM__n120) );
  BUFx2_ASAP7_75t_R EX_MEM___U156 ( .A(EX_ALU_result[22]), .Y(EX_MEM__n235) );
  INVx1_ASAP7_75t_R EX_MEM___U157 ( .A(EX_MEM__n235), .Y(EX_MEM__n121) );
  BUFx2_ASAP7_75t_R EX_MEM___U158 ( .A(EX_ALU_result[20]), .Y(EX_MEM__n237) );
  INVx1_ASAP7_75t_R EX_MEM___U159 ( .A(EX_MEM__n237), .Y(EX_MEM__n122) );
  BUFx2_ASAP7_75t_R EX_MEM___U160 ( .A(EX_ALU_result[16]), .Y(EX_MEM__n241) );
  INVx1_ASAP7_75t_R EX_MEM___U161 ( .A(EX_MEM__n241), .Y(EX_MEM__n123) );
  BUFx2_ASAP7_75t_R EX_MEM___U162 ( .A(EX_ALU_result[15]), .Y(EX_MEM__n242) );
  INVx1_ASAP7_75t_R EX_MEM___U163 ( .A(EX_MEM__n242), .Y(EX_MEM__n124) );
  BUFx2_ASAP7_75t_R EX_MEM___U164 ( .A(EX_ALU_result[13]), .Y(EX_MEM__n244) );
  INVx1_ASAP7_75t_R EX_MEM___U165 ( .A(EX_MEM__n244), .Y(EX_MEM__n125) );
  BUFx2_ASAP7_75t_R EX_MEM___U166 ( .A(EX_ALU_result[2]), .Y(EX_MEM__n255) );
  INVx1_ASAP7_75t_R EX_MEM___U167 ( .A(EX_MEM__n255), .Y(EX_MEM__n126) );
  BUFx2_ASAP7_75t_R EX_MEM___U168 ( .A(ID_EX_RegWrite), .Y(EX_MEM__n272) );
  INVx1_ASAP7_75t_R EX_MEM___U169 ( .A(EX_MEM__n272), .Y(EX_MEM__n127) );
  BUFx2_ASAP7_75t_R EX_MEM___U170 ( .A(ID_EX_MemRead), .Y(EX_MEM__n278) );
  INVx1_ASAP7_75t_R EX_MEM___U171 ( .A(EX_MEM__n278), .Y(EX_MEM__n128) );
  BUFx2_ASAP7_75t_R EX_MEM___U172 ( .A(EX_ALU_result[31]), .Y(EX_MEM__n226) );
  INVx1_ASAP7_75t_R EX_MEM___U173 ( .A(EX_MEM__n226), .Y(EX_MEM__n129) );
  BUFx2_ASAP7_75t_R EX_MEM___U174 ( .A(EX_ALU_result[6]), .Y(EX_MEM__n251) );
  INVx1_ASAP7_75t_R EX_MEM___U175 ( .A(EX_MEM__n251), .Y(EX_MEM__n130) );
  BUFx2_ASAP7_75t_R EX_MEM___U176 ( .A(EX_ALU_result[4]), .Y(EX_MEM__n253) );
  INVx1_ASAP7_75t_R EX_MEM___U177 ( .A(EX_MEM__n253), .Y(EX_MEM__n131) );
  INVx1_ASAP7_75t_R EX_MEM___U178 ( .A(EX_read_reg_data_2[4]), .Y(EX_MEM__n132) );
  BUFx12f_ASAP7_75t_R EX_MEM___U179 ( .A(EX_MEM__n32), .Y(EX_MEM_rd[2]) );
  BUFx3_ASAP7_75t_R EX_MEM___U180 ( .A(EX_MEM__n136), .Y(EX_MEM__n135) );
  BUFx2_ASAP7_75t_R EX_MEM___U181 ( .A(EX_MEM__n285), .Y(EX_MEM__n136) );
  BUFx3_ASAP7_75t_R EX_MEM___U182 ( .A(EX_MEM__n138), .Y(EX_MEM__n137) );
  BUFx2_ASAP7_75t_R EX_MEM___U183 ( .A(EX_MEM__n287), .Y(EX_MEM__n138) );
  BUFx3_ASAP7_75t_R EX_MEM___U184 ( .A(EX_MEM__n140), .Y(EX_MEM__n139) );
  BUFx2_ASAP7_75t_R EX_MEM___U185 ( .A(EX_MEM__n291), .Y(EX_MEM__n140) );
  BUFx3_ASAP7_75t_R EX_MEM___U186 ( .A(EX_MEM__n142), .Y(EX_MEM__n141) );
  BUFx2_ASAP7_75t_R EX_MEM___U187 ( .A(EX_MEM__n296), .Y(EX_MEM__n142) );
  BUFx3_ASAP7_75t_R EX_MEM___U188 ( .A(EX_MEM__n144), .Y(EX_MEM__n143) );
  BUFx2_ASAP7_75t_R EX_MEM___U189 ( .A(EX_MEM__n301), .Y(EX_MEM__n144) );
  BUFx3_ASAP7_75t_R EX_MEM___U190 ( .A(EX_MEM__n147), .Y(EX_MEM__n146) );
  BUFx2_ASAP7_75t_R EX_MEM___U191 ( .A(EX_MEM__n303), .Y(EX_MEM__n147) );
  BUFx3_ASAP7_75t_R EX_MEM___U192 ( .A(EX_MEM__n149), .Y(EX_MEM__n148) );
  BUFx2_ASAP7_75t_R EX_MEM___U193 ( .A(EX_MEM__n306), .Y(EX_MEM__n149) );
  BUFx3_ASAP7_75t_R EX_MEM___U194 ( .A(EX_MEM__n151), .Y(EX_MEM__n150) );
  BUFx2_ASAP7_75t_R EX_MEM___U195 ( .A(EX_MEM__n307), .Y(EX_MEM__n151) );
  BUFx6f_ASAP7_75t_R EX_MEM___U196 ( .A(EX_MEM__n153), .Y(EX_MEM_ALU_result[29]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U197 ( .A(EX_MEM__n86), .Y(EX_MEM__n153) );
  BUFx6f_ASAP7_75t_R EX_MEM___U198 ( .A(EX_MEM__n155), .Y(EX_MEM_ALU_result[25]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U199 ( .A(EX_MEM__n55), .Y(EX_MEM__n155) );
  BUFx6f_ASAP7_75t_R EX_MEM___U200 ( .A(EX_MEM__n157), .Y(EX_MEM_ALU_result[21]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U201 ( .A(EX_MEM__n57), .Y(EX_MEM__n157) );
  BUFx6f_ASAP7_75t_R EX_MEM___U202 ( .A(EX_MEM__n159), .Y(EX_MEM_ALU_result[17]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U203 ( .A(EX_MEM__n96), .Y(EX_MEM__n159) );
  BUFx6f_ASAP7_75t_R EX_MEM___U204 ( .A(EX_MEM__n161), .Y(EX_MEM_ALU_result[10]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U205 ( .A(EX_MEM__n106), .Y(EX_MEM__n161) );
  BUFx6f_ASAP7_75t_R EX_MEM___U206 ( .A(EX_MEM__n163), .Y(EX_MEM_ALU_result[5]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U207 ( .A(EX_MEM__n63), .Y(EX_MEM__n163) );
  BUFx6f_ASAP7_75t_R EX_MEM___U208 ( .A(EX_MEM__n165), .Y(EX_MEM_ALU_result[31]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U209 ( .A(EX_MEM__n51), .Y(EX_MEM__n165) );
  BUFx6f_ASAP7_75t_R EX_MEM___U210 ( .A(EX_MEM__n167), .Y(EX_MEM_ALU_result[30]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U211 ( .A(EX_MEM__n135), .Y(EX_MEM__n167) );
  BUFx6f_ASAP7_75t_R EX_MEM___U212 ( .A(EX_MEM__n169), .Y(EX_MEM_ALU_result[28]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U213 ( .A(EX_MEM__n137), .Y(EX_MEM__n169) );
  BUFx6f_ASAP7_75t_R EX_MEM___U214 ( .A(EX_MEM__n171), .Y(EX_MEM_ALU_result[27]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U215 ( .A(EX_MEM__n88), .Y(EX_MEM__n171) );
  BUFx6f_ASAP7_75t_R EX_MEM___U216 ( .A(EX_MEM__n173), .Y(EX_MEM_ALU_result[26]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U217 ( .A(EX_MEM__n53), .Y(EX_MEM__n173) );
  BUFx6f_ASAP7_75t_R EX_MEM___U218 ( .A(EX_MEM__n175), .Y(EX_MEM_ALU_result[24]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U219 ( .A(EX_MEM__n139), .Y(EX_MEM__n175) );
  BUFx6f_ASAP7_75t_R EX_MEM___U220 ( .A(EX_MEM__n177), .Y(EX_MEM_ALU_result[23]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U221 ( .A(EX_MEM__n90), .Y(EX_MEM__n177) );
  BUFx6f_ASAP7_75t_R EX_MEM___U222 ( .A(EX_MEM__n179), .Y(EX_MEM_ALU_result[22]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U223 ( .A(EX_MEM__n92), .Y(EX_MEM__n179) );
  BUFx6f_ASAP7_75t_R EX_MEM___U224 ( .A(EX_MEM__n181), .Y(EX_MEM_ALU_result[20]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U225 ( .A(EX_MEM__n94), .Y(EX_MEM__n181) );
  BUFx6f_ASAP7_75t_R EX_MEM___U226 ( .A(EX_MEM__n183), .Y(EX_MEM_ALU_result[19]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U227 ( .A(EX_MEM__n141), .Y(EX_MEM__n183) );
  BUFx6f_ASAP7_75t_R EX_MEM___U228 ( .A(EX_MEM__n185), .Y(EX_MEM_ALU_result[18]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U229 ( .A(EX_MEM__n59), .Y(EX_MEM__n185) );
  BUFx6f_ASAP7_75t_R EX_MEM___U230 ( .A(EX_MEM__n187), .Y(EX_MEM_ALU_result[16]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U231 ( .A(EX_MEM__n98), .Y(EX_MEM__n187) );
  BUFx6f_ASAP7_75t_R EX_MEM___U232 ( .A(EX_MEM__n189), .Y(EX_MEM_ALU_result[15]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U233 ( .A(EX_MEM__n100), .Y(EX_MEM__n189) );
  BUFx6f_ASAP7_75t_R EX_MEM___U234 ( .A(EX_MEM__n191), .Y(EX_MEM_ALU_result[14]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U235 ( .A(EX_MEM__n143), .Y(EX_MEM__n191) );
  BUFx6f_ASAP7_75t_R EX_MEM___U236 ( .A(EX_MEM__n193), .Y(EX_MEM_ALU_result[13]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U237 ( .A(EX_MEM__n102), .Y(EX_MEM__n193) );
  BUFx6f_ASAP7_75t_R EX_MEM___U238 ( .A(EX_MEM__n195), .Y(EX_MEM_ALU_result[12]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U239 ( .A(EX_MEM__n146), .Y(EX_MEM__n195) );
  BUFx6f_ASAP7_75t_R EX_MEM___U240 ( .A(EX_MEM__n197), .Y(EX_MEM_ALU_result[11]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U241 ( .A(EX_MEM__n104), .Y(EX_MEM__n197) );
  BUFx6f_ASAP7_75t_R EX_MEM___U242 ( .A(EX_MEM__n199), .Y(EX_MEM_ALU_result[9]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U243 ( .A(EX_MEM__n148), .Y(EX_MEM__n199) );
  BUFx6f_ASAP7_75t_R EX_MEM___U244 ( .A(EX_MEM__n201), .Y(EX_MEM_ALU_result[8]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U245 ( .A(EX_MEM__n150), .Y(EX_MEM__n201) );
  BUFx6f_ASAP7_75t_R EX_MEM___U246 ( .A(EX_MEM__n203), .Y(EX_MEM_ALU_result[7]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U247 ( .A(EX_MEM__n61), .Y(EX_MEM__n203) );
  BUFx6f_ASAP7_75t_R EX_MEM___U248 ( .A(EX_MEM__n205), .Y(EX_MEM_ALU_result[6]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U249 ( .A(EX_MEM__n108), .Y(EX_MEM__n205) );
  BUFx6f_ASAP7_75t_R EX_MEM___U250 ( .A(EX_MEM__n207), .Y(EX_MEM_ALU_result[4]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U251 ( .A(EX_MEM__n65), .Y(EX_MEM__n207) );
  BUFx6f_ASAP7_75t_R EX_MEM___U252 ( .A(EX_MEM__n209), .Y(EX_MEM_ALU_result[3]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U253 ( .A(EX_MEM__n110), .Y(EX_MEM__n209) );
  BUFx6f_ASAP7_75t_R EX_MEM___U254 ( .A(EX_MEM__n211), .Y(EX_MEM_ALU_result[2]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U255 ( .A(EX_MEM__n67), .Y(EX_MEM__n211) );
  BUFx6f_ASAP7_75t_R EX_MEM___U256 ( .A(EX_MEM__n213), .Y(EX_MEM_ALU_result[1]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U257 ( .A(EX_MEM__n112), .Y(EX_MEM__n213) );
  BUFx6f_ASAP7_75t_R EX_MEM___U258 ( .A(EX_MEM__n215), .Y(EX_MEM_ALU_result[0]) );
  BUFx4f_ASAP7_75t_R EX_MEM___U259 ( .A(EX_MEM__n114), .Y(EX_MEM__n215) );
  BUFx4f_ASAP7_75t_R EX_MEM___U260 ( .A(EX_MEM__n26), .Y(EX_MEM__n217) );
  BUFx4f_ASAP7_75t_R EX_MEM___U261 ( .A(EX_MEM__n17), .Y(EX_MEM__n219) );
  BUFx4f_ASAP7_75t_R EX_MEM___U262 ( .A(EX_MEM__n30), .Y(EX_MEM__n221) );
  BUFx12f_ASAP7_75t_R EX_MEM___U263 ( .A(EX_MEM__n223), .Y(EX_MEM_rd[1]) );
  BUFx12f_ASAP7_75t_R EX_MEM___U264 ( .A(EX_MEM__n34), .Y(EX_MEM__n223) );
  BUFx4f_ASAP7_75t_R EX_MEM___U265 ( .A(EX_MEM__n21), .Y(EX_MEM__n225) );
  INVx1_ASAP7_75t_R EX_MEM___U266 ( .A(ID_EX_rd[0]), .Y(EX_MEM__n277) );
  INVx1_ASAP7_75t_R EX_MEM___U267 ( .A(ID_EX_rd[1]), .Y(EX_MEM__n276) );
  INVx1_ASAP7_75t_R EX_MEM___U268 ( .A(ID_EX_rd[3]), .Y(EX_MEM__n274) );
  INVx1_ASAP7_75t_R EX_MEM___U269 ( .A(ID_EX_rd[4]), .Y(EX_MEM__n273) );
  INVx1_ASAP7_75t_R EX_MEM___U270 ( .A(EX_read_reg_data_2[13]), .Y(EX_MEM__n258) );
  INVx1_ASAP7_75t_R EX_MEM___U271 ( .A(EX_read_reg_data_2[14]), .Y(EX_MEM__n259) );
  INVx1_ASAP7_75t_R EX_MEM___U272 ( .A(EX_read_reg_data_2[17]), .Y(EX_MEM__n260) );
  INVx1_ASAP7_75t_R EX_MEM___U273 ( .A(EX_read_reg_data_2[22]), .Y(EX_MEM__n264) );
  INVx1_ASAP7_75t_R EX_MEM___U274 ( .A(EX_read_reg_data_2[31]), .Y(EX_MEM__n268) );
  INVx1_ASAP7_75t_R EX_MEM___U275 ( .A(EX_ALU_result[3]), .Y(EX_MEM__n254) );
  INVx1_ASAP7_75t_R EX_MEM___U276 ( .A(EX_ALU_result[7]), .Y(EX_MEM__n250) );
  INVx1_ASAP7_75t_R EX_MEM___U277 ( .A(EX_ALU_result[24]), .Y(EX_MEM__n233) );
  INVx1_ASAP7_75t_R EX_MEM___U278 ( .A(EX_ALU_result[25]), .Y(EX_MEM__n232) );
  INVx1_ASAP7_75t_R EX_MEM___U279 ( .A(EX_ALU_result[26]), .Y(EX_MEM__n231) );
  INVx1_ASAP7_75t_R EX_MEM___U280 ( .A(EX_ALU_result[27]), .Y(EX_MEM__n230) );
  INVx1_ASAP7_75t_R EX_MEM___U281 ( .A(ID_EX_MemWrite), .Y(EX_MEM__n280) );
  INVx1_ASAP7_75t_R EX_MEM___U282 ( .A(ID_EX_MemToReg), .Y(EX_MEM__n279) );

 BUFx12f_ASAP7_75t_R MEM___U1 ( .A(data_i[26]), .Y(MEM_mem_data[26]) );
  BUFx12f_ASAP7_75t_R MEM___U2 ( .A(data_i[24]), .Y(MEM_mem_data[24]) );
  BUFx12f_ASAP7_75t_R MEM___U3 ( .A(data_i[31]), .Y(MEM_mem_data[31]) );
  BUFx12f_ASAP7_75t_R MEM___U4 ( .A(data_i[23]), .Y(MEM_mem_data[23]) );
  BUFx12f_ASAP7_75t_R MEM___U5 ( .A(data_i[22]), .Y(MEM_mem_data[22]) );
  BUFx12f_ASAP7_75t_R MEM___U6 ( .A(data_i[20]), .Y(MEM_mem_data[20]) );
  BUFx12f_ASAP7_75t_R MEM___U7 ( .A(data_i[18]), .Y(MEM_mem_data[18]) );
  BUFx12f_ASAP7_75t_R MEM___U8 ( .A(data_i[16]), .Y(MEM_mem_data[16]) );
  BUFx12f_ASAP7_75t_R MEM___U9 ( .A(data_i[15]), .Y(MEM_mem_data[15]) );
  BUFx12f_ASAP7_75t_R MEM___U10 ( .A(data_i[13]), .Y(MEM_mem_data[13]) );
  BUFx12f_ASAP7_75t_R MEM___U11 ( .A(data_i[9]), .Y(MEM_mem_data[9]) );
  BUFx12f_ASAP7_75t_R MEM___U12 ( .A(data_i[8]), .Y(MEM_mem_data[8]) );
  BUFx12f_ASAP7_75t_R MEM___U13 ( .A(data_i[6]), .Y(MEM_mem_data[6]) );
  BUFx12f_ASAP7_75t_R MEM___U14 ( .A(data_i[4]), .Y(MEM_mem_data[4]) );
  BUFx12f_ASAP7_75t_R MEM___U15 ( .A(data_i[2]), .Y(MEM_mem_data[2]) );
  BUFx12f_ASAP7_75t_R MEM___U16 ( .A(data_i[0]), .Y(MEM_mem_data[0]) );
  HB1xp67_ASAP7_75t_R MEM___U17 ( .A(EX_MEM_ALU_result[29]), .Y(data_addr_o[29]) );
  HB1xp67_ASAP7_75t_R MEM___U18 ( .A(EX_MEM_ALU_result[25]), .Y(data_addr_o[25]) );
  HB1xp67_ASAP7_75t_R MEM___U19 ( .A(EX_MEM_ALU_result[21]), .Y(data_addr_o[21]) );
  HB1xp67_ASAP7_75t_R MEM___U20 ( .A(EX_MEM_ALU_result[17]), .Y(data_addr_o[17]) );
  HB1xp67_ASAP7_75t_R MEM___U21 ( .A(EX_MEM_ALU_result[10]), .Y(data_addr_o[10]) );
  HB1xp67_ASAP7_75t_R MEM___U22 ( .A(EX_MEM_ALU_result[5]), .Y(data_addr_o[5]) );
  BUFx12f_ASAP7_75t_R MEM___U23 ( .A(data_i[30]), .Y(MEM_mem_data[30]) );
  BUFx12f_ASAP7_75t_R MEM___U24 ( .A(data_i[29]), .Y(MEM_mem_data[29]) );
  BUFx12f_ASAP7_75t_R MEM___U25 ( .A(data_i[28]), .Y(MEM_mem_data[28]) );
  BUFx12f_ASAP7_75t_R MEM___U26 ( .A(data_i[27]), .Y(MEM_mem_data[27]) );
  BUFx12f_ASAP7_75t_R MEM___U27 ( .A(data_i[25]), .Y(MEM_mem_data[25]) );
  BUFx12f_ASAP7_75t_R MEM___U28 ( .A(data_i[21]), .Y(MEM_mem_data[21]) );
  BUFx12f_ASAP7_75t_R MEM___U29 ( .A(data_i[19]), .Y(MEM_mem_data[19]) );
  BUFx12f_ASAP7_75t_R MEM___U30 ( .A(data_i[17]), .Y(MEM_mem_data[17]) );
  BUFx12f_ASAP7_75t_R MEM___U31 ( .A(data_i[14]), .Y(MEM_mem_data[14]) );
  BUFx12f_ASAP7_75t_R MEM___U32 ( .A(data_i[12]), .Y(MEM_mem_data[12]) );
  BUFx12f_ASAP7_75t_R MEM___U33 ( .A(data_i[11]), .Y(MEM_mem_data[11]) );
  BUFx12f_ASAP7_75t_R MEM___U34 ( .A(data_i[10]), .Y(MEM_mem_data[10]) );
  BUFx12f_ASAP7_75t_R MEM___U35 ( .A(data_i[7]), .Y(MEM_mem_data[7]) );
  BUFx12f_ASAP7_75t_R MEM___U36 ( .A(data_i[5]), .Y(MEM_mem_data[5]) );
  BUFx12f_ASAP7_75t_R MEM___U37 ( .A(data_i[3]), .Y(MEM_mem_data[3]) );
  BUFx12f_ASAP7_75t_R MEM___U38 ( .A(data_i[1]), .Y(MEM_mem_data[1]) );
  HB1xp67_ASAP7_75t_R MEM___U39 ( .A(n74), .Y(data_o[30]) );
  HB1xp67_ASAP7_75t_R MEM___U40 ( .A(n75), .Y(data_o[28]) );
  HB1xp67_ASAP7_75t_R MEM___U41 ( .A(n76), .Y(data_o[19]) );
  HB1xp67_ASAP7_75t_R MEM___U42 ( .A(n94), .Y(data_we_o) );
  HB1xp67_ASAP7_75t_R MEM___U43 ( .A(n95), .Y(data_o[31]) );
  HB1xp67_ASAP7_75t_R MEM___U44 ( .A(n96), .Y(data_o[29]) );
  HB1xp67_ASAP7_75t_R MEM___U45 ( .A(n97), .Y(data_o[27]) );
  HB1xp67_ASAP7_75t_R MEM___U46 ( .A(n98), .Y(data_o[26]) );
  HB1xp67_ASAP7_75t_R MEM___U47 ( .A(n99), .Y(data_o[25]) );
  HB1xp67_ASAP7_75t_R MEM___U48 ( .A(n100), .Y(data_o[24]) );
  HB1xp67_ASAP7_75t_R MEM___U49 ( .A(n101), .Y(data_o[23]) );
  HB1xp67_ASAP7_75t_R MEM___U50 ( .A(n102), .Y(data_o[22]) );
  HB1xp67_ASAP7_75t_R MEM___U51 ( .A(n103), .Y(data_o[21]) );
  HB1xp67_ASAP7_75t_R MEM___U52 ( .A(n104), .Y(data_o[20]) );
  HB1xp67_ASAP7_75t_R MEM___U53 ( .A(n105), .Y(data_o[18]) );
  HB1xp67_ASAP7_75t_R MEM___U54 ( .A(n106), .Y(data_o[17]) );
  HB1xp67_ASAP7_75t_R MEM___U55 ( .A(n107), .Y(data_o[16]) );
  HB1xp67_ASAP7_75t_R MEM___U56 ( .A(EX_MEM_ALU_result[31]), .Y(data_addr_o[31]) );
  HB1xp67_ASAP7_75t_R MEM___U57 ( .A(EX_MEM_ALU_result[30]), .Y(data_addr_o[30]) );
  HB1xp67_ASAP7_75t_R MEM___U58 ( .A(EX_MEM_ALU_result[28]), .Y(data_addr_o[28]) );
  HB1xp67_ASAP7_75t_R MEM___U59 ( .A(EX_MEM_ALU_result[27]), .Y(data_addr_o[27]) );
  HB1xp67_ASAP7_75t_R MEM___U60 ( .A(EX_MEM_ALU_result[26]), .Y(data_addr_o[26]) );
  HB1xp67_ASAP7_75t_R MEM___U61 ( .A(EX_MEM_ALU_result[24]), .Y(data_addr_o[24]) );
  HB1xp67_ASAP7_75t_R MEM___U62 ( .A(EX_MEM_ALU_result[23]), .Y(data_addr_o[23]) );
  HB1xp67_ASAP7_75t_R MEM___U63 ( .A(EX_MEM_ALU_result[22]), .Y(data_addr_o[22]) );
  HB1xp67_ASAP7_75t_R MEM___U64 ( .A(EX_MEM_ALU_result[20]), .Y(data_addr_o[20]) );
  HB1xp67_ASAP7_75t_R MEM___U65 ( .A(EX_MEM_ALU_result[19]), .Y(data_addr_o[19]) );
  HB1xp67_ASAP7_75t_R MEM___U66 ( .A(EX_MEM_ALU_result[18]), .Y(data_addr_o[18]) );
  HB1xp67_ASAP7_75t_R MEM___U67 ( .A(EX_MEM_ALU_result[16]), .Y(data_addr_o[16]) );
  HB1xp67_ASAP7_75t_R MEM___U68 ( .A(EX_MEM_ALU_result[15]), .Y(data_addr_o[15]) );
  HB1xp67_ASAP7_75t_R MEM___U69 ( .A(EX_MEM_ALU_result[14]), .Y(data_addr_o[14]) );
  HB1xp67_ASAP7_75t_R MEM___U70 ( .A(EX_MEM_ALU_result[13]), .Y(data_addr_o[13]) );
  HB1xp67_ASAP7_75t_R MEM___U71 ( .A(EX_MEM_ALU_result[12]), .Y(data_addr_o[12]) );
  HB1xp67_ASAP7_75t_R MEM___U72 ( .A(EX_MEM_ALU_result[11]), .Y(data_addr_o[11]) );
  HB1xp67_ASAP7_75t_R MEM___U73 ( .A(EX_MEM_ALU_result[9]), .Y(data_addr_o[9]) );
  HB1xp67_ASAP7_75t_R MEM___U74 ( .A(EX_MEM_ALU_result[8]), .Y(data_addr_o[8]) );
  HB1xp67_ASAP7_75t_R MEM___U75 ( .A(EX_MEM_ALU_result[7]), .Y(data_addr_o[7]) );
  HB1xp67_ASAP7_75t_R MEM___U76 ( .A(EX_MEM_ALU_result[6]), .Y(data_addr_o[6]) );
  HB1xp67_ASAP7_75t_R MEM___U77 ( .A(EX_MEM_ALU_result[4]), .Y(data_addr_o[4]) );
  HB1xp67_ASAP7_75t_R MEM___U78 ( .A(EX_MEM_ALU_result[3]), .Y(data_addr_o[3]) );
  HB1xp67_ASAP7_75t_R MEM___U79 ( .A(EX_MEM_ALU_result[2]), .Y(data_addr_o[2]) );
  HB1xp67_ASAP7_75t_R MEM___U80 ( .A(EX_MEM_ALU_result[1]), .Y(data_addr_o[1]) );
  HB1xp67_ASAP7_75t_R MEM___U81 ( .A(EX_MEM_ALU_result[0]), .Y(data_addr_o[0]) );
  HB1xp67_ASAP7_75t_R MEM___U82 ( .A(n82), .Y(data_o[15]) );
  HB1xp67_ASAP7_75t_R MEM___U83 ( .A(n77), .Y(data_o[14]) );
  HB1xp67_ASAP7_75t_R MEM___U84 ( .A(n83), .Y(data_o[13]) );
  HB1xp67_ASAP7_75t_R MEM___U85 ( .A(n84), .Y(data_o[12]) );
  HB1xp67_ASAP7_75t_R MEM___U86 ( .A(n78), .Y(data_o[11]) );
  HB1xp67_ASAP7_75t_R MEM___U87 ( .A(n85), .Y(data_o[10]) );
  HB1xp67_ASAP7_75t_R MEM___U88 ( .A(n86), .Y(data_o[9]) );
  HB1xp67_ASAP7_75t_R MEM___U89 ( .A(n87), .Y(data_o[8]) );
  HB1xp67_ASAP7_75t_R MEM___U90 ( .A(n88), .Y(data_o[7]) );
  HB1xp67_ASAP7_75t_R MEM___U91 ( .A(n89), .Y(data_o[6]) );
  HB1xp67_ASAP7_75t_R MEM___U92 ( .A(n90), .Y(data_o[5]) );
  HB1xp67_ASAP7_75t_R MEM___U93 ( .A(n91), .Y(data_o[4]) );
  HB1xp67_ASAP7_75t_R MEM___U94 ( .A(n79), .Y(data_o[3]) );
  HB1xp67_ASAP7_75t_R MEM___U95 ( .A(n92), .Y(data_o[2]) );
  HB1xp67_ASAP7_75t_R MEM___U96 ( .A(n80), .Y(data_o[1]) );
  HB1xp67_ASAP7_75t_R MEM___U97 ( .A(n93), .Y(data_o[0]) );

   DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_31_ ( .D(MEM_WB__n253), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n286) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_30_ ( .D(MEM_WB__n254), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n287) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_29_ ( .D(MEM_WB__n255), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n288) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_28_ ( .D(MEM_WB__n256), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n289) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_27_ ( .D(MEM_WB__n257), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n290) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_26_ ( .D(MEM_WB__n258), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n291) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_25_ ( .D(MEM_WB__n259), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(mem_data_out[25]) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_24_ ( .D(MEM_WB__n260), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(mem_data_out[24]) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_23_ ( .D(MEM_WB__n261), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n292) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_22_ ( .D(MEM_WB__n262), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n293) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_21_ ( .D(MEM_WB__n263), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n294) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_20_ ( .D(MEM_WB__n264), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n295) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_19_ ( .D(MEM_WB__n265), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n296) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_18_ ( .D(MEM_WB__n266), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n297) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_17_ ( .D(MEM_WB__n267), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n298) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_16_ ( .D(MEM_WB__n268), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(mem_data_out[16]) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_15_ ( .D(MEM_WB__n269), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n299) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_14_ ( .D(MEM_WB__n270), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n300) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_13_ ( .D(MEM_WB__n271), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n301) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_12_ ( .D(MEM_WB__n272), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n302) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_11_ ( .D(MEM_WB__n273), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n303) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_10_ ( .D(MEM_WB__n274), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n304) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_9_ ( .D(MEM_WB__n275), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n305) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_8_ ( .D(MEM_WB__n276), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n306) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_7_ ( .D(MEM_WB__n277), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n307) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_6_ ( .D(MEM_WB__n278), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n308) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_5_ ( .D(MEM_WB__n279), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n309) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_4_ ( .D(MEM_WB__n280), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(mem_data_out[4]) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_3_ ( .D(MEM_WB__n281), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n310) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_2_ ( .D(MEM_WB__n282), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n311) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_1_ ( .D(MEM_WB__n283), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n312) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___mem_data_out_reg_0_ ( .D(MEM_WB__n284), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n313) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___rd_out_reg_3_ ( .D(MEM_WB__n155), .CLK(clk), .SETN(MEM_WB__n143), 
        .RESETN(MEM_WB__n212), .QN(MEM_WB_rd[3]) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___rd_out_reg_2_ ( .D(MEM_WB__n156), .CLK(clk), .SETN(MEM_WB__n143), 
        .RESETN(MEM_WB__n212), .QN(MEM_WB_rd[2]) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_31_ ( .D(MEM_WB__n219), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n314) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_30_ ( .D(MEM_WB__n220), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n315) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_29_ ( .D(MEM_WB__n184), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n316) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_28_ ( .D(MEM_WB__n222), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n317) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_27_ ( .D(MEM_WB__n61), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n318) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_26_ ( .D(MEM_WB__n224), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n319) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_25_ ( .D(MEM_WB__n185), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n320) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_24_ ( .D(MEM_WB__n28), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n321) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_23_ ( .D(MEM_WB__n37), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n322) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_22_ ( .D(MEM_WB__n228), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n323) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_21_ ( .D(MEM_WB__n186), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n324) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_20_ ( .D(MEM_WB__n29), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n325) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_19_ ( .D(MEM_WB__n231), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n326) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_18_ ( .D(MEM_WB__n24), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n327) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_17_ ( .D(MEM_WB__n187), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n328) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_16_ ( .D(MEM_WB__n30), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n329) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_15_ ( .D(MEM_WB__n235), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n330) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_14_ ( .D(MEM_WB__n236), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n331) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_13_ ( .D(MEM_WB__n237), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n332) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_12_ ( .D(MEM_WB__n238), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n333) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_11_ ( .D(MEM_WB__n239), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n334) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_10_ ( .D(MEM_WB__n188), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n335) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_9_ ( .D(MEM_WB__n31), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n336) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_8_ ( .D(MEM_WB__n242), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n337) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_7_ ( .D(MEM_WB__n243), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n338) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_6_ ( .D(MEM_WB__n244), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n339) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_5_ ( .D(MEM_WB__n189), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n340) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_4_ ( .D(MEM_WB__n246), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n341) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_3_ ( .D(MEM_WB__n247), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n342) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_2_ ( .D(MEM_WB__n23), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n343) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_1_ ( .D(MEM_WB__n249), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n344) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___ALU_result_out_reg_0_ ( .D(MEM_WB__n250), .CLK(clk), .SETN(
        n143), .RESETN(MEM_WB__n212), .QN(MEM_WB__n345) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___MemRead_out_reg ( .D(MEM_WB__n251), .CLK(clk), .SETN(MEM_WB__n143), 
        .RESETN(MEM_WB__n212), .QN(MEM_WB_MemRead) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___MemtoReg_out_reg ( .D(MEM_WB__n252), .CLK(clk), .SETN(MEM_WB__n143), 
        .RESETN(MEM_WB__n212), .QN(MEM_WB_MemtoReg) );
  CKINVDCx10_ASAP7_75t_R MEM_WB___U145 ( .A(rst), .Y(MEM_WB__n143) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___RegWrite_out_reg ( .D(MEM_WB__n218), .CLK(clk), .SETN(MEM_WB__n143), 
        .RESETN(MEM_WB__n212), .QN(MEM_WB__n285) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___rd_out_reg_1_ ( .D(MEM_WB__n22), .CLK(clk), .SETN(MEM_WB__n143), 
        .RESETN(MEM_WB__n212), .QN(MEM_WB_rd[1]) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___rd_out_reg_0_ ( .D(MEM_WB__n122), .CLK(clk), .SETN(MEM_WB__n143), 
        .RESETN(MEM_WB__n212), .QN(MEM_WB__n346) );
  DFFASRHQNx1_ASAP7_75t_R MEM_WB___rd_out_reg_4_ ( .D(MEM_WB__n157), .CLK(clk), .SETN(MEM_WB__n143), 
        .RESETN(MEM_WB__n212), .QN(MEM_WB_rd[4]) );
  TIEHIx1_ASAP7_75t_R MEM_WB___U3 ( .H(MEM_WB__n212) );
  BUFx2_ASAP7_75t_R MEM_WB___U4 ( .A(MEM_WB__n144), .Y(mem_data_out[1]) );
  BUFx3_ASAP7_75t_R MEM_WB___U5 ( .A(MEM_WB__n59), .Y(MEM_WB_ALU_result[9]) );
  BUFx3_ASAP7_75t_R MEM_WB___U6 ( .A(MEM_WB__n207), .Y(mem_data_out[9]) );
  BUFx2_ASAP7_75t_R MEM_WB___U7 ( .A(MEM_WB__n63), .Y(MEM_WB__n201) );
  HB1xp67_ASAP7_75t_R MEM_WB___U8 ( .A(MEM_WB__n32), .Y(MEM_WB__n199) );
  HB1xp67_ASAP7_75t_R MEM_WB___U9 ( .A(MEM_WB__n199), .Y(mem_data_out[13]) );
  HB1xp67_ASAP7_75t_R MEM_WB___U10 ( .A(MEM_WB__n306), .Y(MEM_WB__n63) );
  BUFx12f_ASAP7_75t_R MEM_WB___U11 ( .A(MEM_WB__n211), .Y(mem_data_out[0]) );
  BUFx6f_ASAP7_75t_R MEM_WB___U12 ( .A(MEM_WB__n126), .Y(MEM_WB__n211) );
  BUFx6f_ASAP7_75t_R MEM_WB___U13 ( .A(MEM_WB__n167), .Y(MEM_WB_ALU_result[13]) );
  HB1xp67_ASAP7_75t_R MEM_WB___U14 ( .A(MEM_WB__n124), .Y(MEM_WB__n32) );
  BUFx3_ASAP7_75t_R MEM_WB___U15 ( .A(MEM_WB__n177), .Y(MEM_WB_ALU_result[3]) );
  BUFx3_ASAP7_75t_R MEM_WB___U16 ( .A(MEM_WB__n140), .Y(mem_data_out[3]) );
  BUFx3_ASAP7_75t_R MEM_WB___U17 ( .A(MEM_WB__n195), .Y(mem_data_out[18]) );
  HB1xp67_ASAP7_75t_R MEM_WB___U18 ( .A(MEM_WB__n35), .Y(MEM_WB__n144) );
  BUFx2_ASAP7_75t_R MEM_WB___U19 ( .A(MEM_WB__n25), .Y(MEM_WB__n195) );
  BUFx6f_ASAP7_75t_R MEM_WB___U20 ( .A(MEM_WB__n193), .Y(mem_data_out[20]) );
  BUFx3_ASAP7_75t_R MEM_WB___U21 ( .A(MEM_WB__n161), .Y(MEM_WB_ALU_result[20]) );
  HB1xp67_ASAP7_75t_R MEM_WB___U22 ( .A(MEM_WB__n112), .Y(MEM_WB__n25) );
  BUFx6f_ASAP7_75t_R MEM_WB___U23 ( .A(MEM_WB__n21), .Y(MEM_WB__n80) );
  BUFx12f_ASAP7_75t_R MEM_WB___U24 ( .A(MEM_WB__n80), .Y(mem_data_out[27]) );
  HB1xp67_ASAP7_75t_R MEM_WB___U25 ( .A(MEM_WB__n297), .Y(MEM_WB__n112) );
  HB1xp67_ASAP7_75t_R MEM_WB___U26 ( .A(MEM_WB__n301), .Y(MEM_WB__n124) );
  BUFx3_ASAP7_75t_R MEM_WB___U27 ( .A(MEM_WB__n138), .Y(mem_data_out[19]) );
  HB1xp67_ASAP7_75t_R MEM_WB___U28 ( .A(MEM_WB__n311), .Y(MEM_WB__n114) );
  BUFx6f_ASAP7_75t_R MEM_WB___U29 ( .A(MEM_WB__n209), .Y(mem_data_out[2]) );
  BUFx3_ASAP7_75t_R MEM_WB___U30 ( .A(MEM_WB__n346), .Y(MEM_WB_rd[0]) );
  HB1xp67_ASAP7_75t_R MEM_WB___U31 ( .A(MEM_WB__n103), .Y(MEM_WB__n159) );
  HB1xp67_ASAP7_75t_R MEM_WB___U32 ( .A(MEM_WB__n323), .Y(MEM_WB__n103) );
  HB1xp67_ASAP7_75t_R MEM_WB___U33 ( .A(MEM_WB__n181), .Y(MEM_WB_ALU_result[1]) );
  HB1xp67_ASAP7_75t_R MEM_WB___U34 ( .A(MEM_WB__n312), .Y(MEM_WB__n35) );
  BUFx3_ASAP7_75t_R MEM_WB___U35 ( .A(MEM_WB__n285), .Y(MEM_WB_RegWrite) );
  HB1xp67_ASAP7_75t_R MEM_WB___U36 ( .A(MEM_WB__n322), .Y(MEM_WB__n11) );
  HB1xp67_ASAP7_75t_R MEM_WB___U37 ( .A(MEM_WB__n292), .Y(MEM_WB__n39) );
  HB1xp67_ASAP7_75t_R MEM_WB___U38 ( .A(MEM_WB__n48), .Y(MEM_WB__n181) );
  HB1xp67_ASAP7_75t_R MEM_WB___U39 ( .A(MEM_WB__n340), .Y(MEM_WB__n101) );
  HB1xp67_ASAP7_75t_R MEM_WB___U40 ( .A(MEM_WB__n344), .Y(MEM_WB__n48) );
  BUFx12f_ASAP7_75t_R MEM_WB___U41 ( .A(MEM_WB__n150), .Y(MEM_WB_ALU_result[25]) );
  BUFx3_ASAP7_75t_R MEM_WB___U42 ( .A(MEM_WB__n169), .Y(MEM_WB_ALU_result[6]) );
  BUFx12f_ASAP7_75t_R MEM_WB___U43 ( .A(MEM_WB__n134), .Y(MEM_WB_ALU_result[5]) );
  BUFx6f_ASAP7_75t_R MEM_WB___U44 ( .A(MEM_WB__n100), .Y(MEM_WB__n134) );
  HB1xp67_ASAP7_75t_R MEM_WB___U45 ( .A(MEM_WB__n303), .Y(MEM_WB__n41) );
  BUFx6f_ASAP7_75t_R MEM_WB___U46 ( .A(MEM_WB__n109), .Y(mem_data_out[11]) );
  HB1xp67_ASAP7_75t_R MEM_WB___U47 ( .A(MEM_WB__n325), .Y(MEM_WB__n115) );
  BUFx2_ASAP7_75t_R MEM_WB___U48 ( .A(MEM_WB__n82), .Y(mem_data_out[17]) );
  HB1xp67_ASAP7_75t_R MEM_WB___U49 ( .A(MEM_WB__MEM_WB__n328), .Y(MEM_WB__n3) );
  HB1xp67_ASAP7_75t_R MEM_WB___U50 ( .A(MEM_WB__n16), .Y(MEM_WB__n82) );
  HB1xp67_ASAP7_75t_R MEM_WB___U51 ( .A(MEM_WB__n298), .Y(MEM_WB__n16) );
  BUFx3_ASAP7_75t_R MEM_WB___U52 ( .A(MEM_WB__n128), .Y(MEM_WB_ALU_result[21]) );
  BUFx6f_ASAP7_75t_R MEM_WB___U53 ( .A(MEM_WB__n132), .Y(MEM_WB_ALU_result[8]) );
  BUFx6f_ASAP7_75t_R MEM_WB___U54 ( .A(MEM_WB__n201), .Y(mem_data_out[8]) );
  BUFx2_ASAP7_75t_R MEM_WB___U55 ( .A(MEM_WB__n316), .Y(MEM_WB__n1) );
  BUFx4f_ASAP7_75t_R MEM_WB___U56 ( .A(MEM_WB__n51), .Y(MEM_WB_ALU_result[29]) );
  BUFx3_ASAP7_75t_R MEM_WB___U57 ( .A(MEM_WB__n1), .Y(MEM_WB__n51) );
  BUFx2_ASAP7_75t_R MEM_WB___U58 ( .A(MEM_WB__n321), .Y(MEM_WB__n2) );
  BUFx4f_ASAP7_75t_R MEM_WB___U59 ( .A(MEM_WB__n68), .Y(MEM_WB_ALU_result[24]) );
  BUFx3_ASAP7_75t_R MEM_WB___U60 ( .A(MEM_WB__n2), .Y(MEM_WB__n68) );
  BUFx4f_ASAP7_75t_R MEM_WB___U61 ( .A(MEM_WB__n55), .Y(MEM_WB_ALU_result[17]) );
  BUFx3_ASAP7_75t_R MEM_WB___U62 ( .A(MEM_WB__n3), .Y(MEM_WB__n55) );
  BUFx2_ASAP7_75t_R MEM_WB___U63 ( .A(MEM_WB__n333), .Y(MEM_WB__n4) );
  BUFx4f_ASAP7_75t_R MEM_WB___U64 ( .A(MEM_WB__n57), .Y(MEM_WB_ALU_result[12]) );
  BUFx3_ASAP7_75t_R MEM_WB___U65 ( .A(MEM_WB__n4), .Y(MEM_WB__n57) );
  BUFx2_ASAP7_75t_R MEM_WB___U66 ( .A(MEM_WB__n336), .Y(MEM_WB__n5) );
  BUFx3_ASAP7_75t_R MEM_WB___U67 ( .A(MEM_WB__n5), .Y(MEM_WB__MEM_WB__n59) );
  BUFx2_ASAP7_75t_R MEM_WB___U68 ( .A(MEM_WB__n304), .Y(MEM_WB__n6) );
  BUFx2_ASAP7_75t_R MEM_WB___U69 ( .A(MEM_WB__n289), .Y(MEM_WB__n7) );
  BUFx2_ASAP7_75t_R MEM_WB___U70 ( .A(MEM_WB__n317), .Y(MEM_WB__n8) );
  BUFx2_ASAP7_75t_R MEM_WB___U71 ( .A(MEM_WB__n318), .Y(MEM_WB__n10) );
  BUFx4f_ASAP7_75t_R MEM_WB___U72 ( .A(MEM_WB__n53), .Y(MEM_WB_ALU_result[27]) );
  BUFx3_ASAP7_75t_R MEM_WB___U73 ( .A(MEM_WB__n10), .Y(MEM_WB__n53) );
  BUFx4f_ASAP7_75t_R MEM_WB___U74 ( .A(MEM_WB__n70), .Y(MEM_WB_ALU_result[23]) );
  BUFx3_ASAP7_75t_R MEM_WB___U75 ( .A(MEM_WB__n11), .Y(MEM_WB__n70) );
  BUFx2_ASAP7_75t_R MEM_WB___U76 ( .A(MEM_WB__n326), .Y(MEM_WB__n12) );
  BUFx4f_ASAP7_75t_R MEM_WB___U77 ( .A(MEM_WB__n72), .Y(MEM_WB_ALU_result[19]) );
  BUFx3_ASAP7_75t_R MEM_WB___U78 ( .A(MEM_WB__n12), .Y(MEM_WB__n72) );
  BUFx2_ASAP7_75t_R MEM_WB___U79 ( .A(MEM_WB__n286), .Y(MEM_WB__n13) );
  BUFx2_ASAP7_75t_R MEM_WB___U80 ( .A(MEM_WB__n287), .Y(MEM_WB__n14) );
  BUFx2_ASAP7_75t_R MEM_WB___U81 ( .A(MEM_WB__n288), .Y(MEM_WB__n15) );
  BUFx2_ASAP7_75t_R MEM_WB___U82 ( .A(MEM_WB__n300), .Y(MEM_WB__n17) );
  BUFx2_ASAP7_75t_R MEM_WB___U83 ( .A(MEM_WB__n302), .Y(MEM_WB__n18) );
  BUFx2_ASAP7_75t_R MEM_WB___U84 ( .A(MEM_WB__n305), .Y(MEM_WB__n19) );
  BUFx2_ASAP7_75t_R MEM_WB___U85 ( .A(MEM_WB__n319), .Y(MEM_WB__n20) );
  BUFx4f_ASAP7_75t_R MEM_WB___U86 ( .A(MEM_WB__n66), .Y(MEM_WB_ALU_result[26]) );
  BUFx3_ASAP7_75t_R MEM_WB___U87 ( .A(MEM_WB__n20), .Y(MEM_WB__n66) );
  BUFx2_ASAP7_75t_R MEM_WB___U88 ( .A(MEM_WB__n290), .Y(MEM_WB__n21) );
  BUFx2_ASAP7_75t_R MEM_WB___U89 ( .A(MEM_WB__n216), .Y(MEM_WB__n22) );
  BUFx2_ASAP7_75t_R MEM_WB___U90 ( .A(MEM_WB__n248), .Y(MEM_WB__n23) );
  BUFx2_ASAP7_75t_R MEM_WB___U91 ( .A(MEM_WB__n232), .Y(MEM_WB__n24) );
  BUFx2_ASAP7_75t_R MEM_WB___U92 ( .A(MEM_WB__n307), .Y(MEM_WB__n26) );
  BUFx2_ASAP7_75t_R MEM_WB___U93 ( .A(MEM_WB__n310), .Y(MEM_WB__n27) );
  BUFx2_ASAP7_75t_R MEM_WB___U94 ( .A(MEM_WB__n226), .Y(MEM_WB__n28) );
  BUFx2_ASAP7_75t_R MEM_WB___U95 ( .A(MEM_WB__n230), .Y(MEM_WB__n29) );
  BUFx2_ASAP7_75t_R MEM_WB___U96 ( .A(MEM_WB__n234), .Y(MEM_WB__n30) );
  BUFx2_ASAP7_75t_R MEM_WB___U97 ( .A(MEM_WB__n241), .Y(MEM_WB__n31) );
  BUFx6f_ASAP7_75t_R MEM_WB___U98 ( .A(MEM_WB__n120), .Y(mem_data_out[5]) );
  BUFx4f_ASAP7_75t_R MEM_WB___U99 ( .A(MEM_WB__n121), .Y(MEM_WB__n120) );
  BUFx2_ASAP7_75t_R MEM_WB___U100 ( .A(MEM_WB__n334), .Y(MEM_WB__n34) );
  BUFx4f_ASAP7_75t_R MEM_WB___U101 ( .A(MEM_WB__n74), .Y(MEM_WB_ALU_result[11]) );
  BUFx3_ASAP7_75t_R MEM_WB___U102 ( .A(MEM_WB__n34), .Y(MEM_WB__n74) );
  BUFx2_ASAP7_75t_R MEM_WB___U103 ( .A(MEM_WB__n338), .Y(MEM_WB__n36) );
  BUFx2_ASAP7_75t_R MEM_WB___U104 ( .A(MEM_WB__n227), .Y(MEM_WB__n37) );
  BUFx2_ASAP7_75t_R MEM_WB___U105 ( .A(MEM_WB__n291), .Y(MEM_WB__n38) );
  BUFx2_ASAP7_75t_R MEM_WB___U106 ( .A(MEM_WB__n296), .Y(MEM_WB__n40) );
  BUFx2_ASAP7_75t_R MEM_WB___U107 ( .A(MEM_WB__n314), .Y(MEM_WB__n42) );
  BUFx2_ASAP7_75t_R MEM_WB___U108 ( .A(MEM_WB__n315), .Y(MEM_WB__n43) );
  BUFx2_ASAP7_75t_R MEM_WB___U109 ( .A(MEM_WB__n331), .Y(MEM_WB__n44) );
  BUFx2_ASAP7_75t_R MEM_WB___U110 ( .A(MEM_WB__n332), .Y(MEM_WB__n45) );
  BUFx2_ASAP7_75t_R MEM_WB___U111 ( .A(MEM_WB__n335), .Y(MEM_WB__n46) );
  BUFx2_ASAP7_75t_R MEM_WB___U112 ( .A(MEM_WB__n342), .Y(MEM_WB__n47) );
  BUFx2_ASAP7_75t_R MEM_WB___U113 ( .A(EX_MEM_rd[3]), .Y(MEM_WB__n49) );
  BUFx2_ASAP7_75t_R MEM_WB___U114 ( .A(MEM_WB__n223), .Y(MEM_WB__n61) );
  BUFx2_ASAP7_75t_R MEM_WB___U115 ( .A(MEM_WB__n293), .Y(MEM_WB__n62) );
  BUFx4f_ASAP7_75t_R MEM_WB___U116 ( .A(MEM_WB__n191), .Y(mem_data_out[22]) );
  BUFx3_ASAP7_75t_R MEM_WB___U117 ( .A(MEM_WB__n62), .Y(MEM_WB__n191) );
  BUFx2_ASAP7_75t_R MEM_WB___U118 ( .A(EX_MEM_rd[0]), .Y(MEM_WB__n64) );
  BUFx4f_ASAP7_75t_R MEM_WB___U119 ( .A(MEM_WB__n76), .Y(mem_data_out[30]) );
  BUFx3_ASAP7_75t_R MEM_WB___U120 ( .A(MEM_WB__n14), .Y(MEM_WB__n76) );
  BUFx4f_ASAP7_75t_R MEM_WB___U121 ( .A(MEM_WB__n78), .Y(mem_data_out[28]) );
  BUFx3_ASAP7_75t_R MEM_WB___U122 ( .A(MEM_WB__n7), .Y(MEM_WB__MEM_WB__n78) );
  BUFx4f_ASAP7_75t_R MEM_WB___U123 ( .A(MEM_WB__n84), .Y(mem_data_out[14]) );
  BUFx3_ASAP7_75t_R MEM_WB___U124 ( .A(MEM_WB__n17), .Y(MEM_WB__n84) );
  BUFx4f_ASAP7_75t_R MEM_WB___U125 ( .A(MEM_WB__n86), .Y(mem_data_out[12]) );
  BUFx3_ASAP7_75t_R MEM_WB___U126 ( .A(MEM_WB__n18), .Y(MEM_WB__n86) );
  BUFx4f_ASAP7_75t_R MEM_WB___U127 ( .A(MEM_WB__n88), .Y(mem_data_out[7]) );
  BUFx3_ASAP7_75t_R MEM_WB___U128 ( .A(MEM_WB__n26), .Y(MEM_WB__n88) );
  BUFx4f_ASAP7_75t_R MEM_WB___U129 ( .A(MEM_WB__n90), .Y(MEM_WB_ALU_result[31]) );
  BUFx3_ASAP7_75t_R MEM_WB___U130 ( .A(MEM_WB__n42), .Y(MEM_WB__n90) );
  BUFx4f_ASAP7_75t_R MEM_WB___U131 ( .A(MEM_WB__n92), .Y(MEM_WB_ALU_result[10]) );
  BUFx3_ASAP7_75t_R MEM_WB___U132 ( .A(MEM_WB__n46), .Y(MEM_WB__n92) );
  BUFx2_ASAP7_75t_R MEM_WB___U133 ( .A(MEM_WB__n295), .Y(MEM_WB__n93) );
  BUFx3_ASAP7_75t_R MEM_WB___U134 ( .A(MEM_WB__n93), .Y(MEM_WB__n193) );
  BUFx3_ASAP7_75t_R MEM_WB___U135 ( .A(MEM_WB__n95), .Y(MEM_WB__n94) );
  BUFx2_ASAP7_75t_R MEM_WB___U136 ( .A(MEM_WB__n324), .Y(MEM_WB__n95) );
  BUFx3_ASAP7_75t_R MEM_WB___U137 ( .A(MEM_WB__n94), .Y(MEM_WB__n128) );
  BUFx2_ASAP7_75t_R MEM_WB___U138 ( .A(MEM_WB__n327), .Y(MEM_WB__n96) );
  BUFx4f_ASAP7_75t_R MEM_WB___U139 ( .A(MEM_WB__n130), .Y(MEM_WB_ALU_result[18]) );
  BUFx3_ASAP7_75t_R MEM_WB___U140 ( .A(MEM_WB__n96), .Y(MEM_WB__n130) );
  BUFx2_ASAP7_75t_R MEM_WB___U141 ( .A(MEM_WB__n329), .Y(MEM_WB__n97) );
  BUFx4f_ASAP7_75t_R MEM_WB___U142 ( .A(MEM_WB__n163), .Y(MEM_WB_ALU_result[16]) );
  BUFx3_ASAP7_75t_R MEM_WB___U143 ( .A(MEM_WB__n97), .Y(MEM_WB__n163) );
  BUFx2_ASAP7_75t_R MEM_WB___U144 ( .A(MEM_WB__n330), .Y(MEM_WB__n98) );
  BUFx4f_ASAP7_75t_R MEM_WB___U146 ( .A(MEM_WB__n164), .Y(MEM_WB_ALU_result[15]) );
  BUFx3_ASAP7_75t_R MEM_WB___U147 ( .A(MEM_WB__n101), .Y(MEM_WB__n100) );
  BUFx2_ASAP7_75t_R MEM_WB___U148 ( .A(MEM_WB__n320), .Y(MEM_WB__n102) );
  BUFx2_ASAP7_75t_R MEM_WB___U149 ( .A(MEM_WB__n341), .Y(MEM_WB__n104) );
  BUFx2_ASAP7_75t_R MEM_WB___U150 ( .A(MEM_WB__n343), .Y(MEM_WB__n105) );
  BUFx2_ASAP7_75t_R MEM_WB___U151 ( .A(EX_MEM_rd[4]), .Y(MEM_WB__n106) );
  BUFx2_ASAP7_75t_R MEM_WB___U152 ( .A(EX_MEM_rd[2]), .Y(MEM_WB__n107) );
  BUFx3_ASAP7_75t_R MEM_WB___U153 ( .A(MEM_WB__n41), .Y(MEM_WB__n109) );
  BUFx4f_ASAP7_75t_R MEM_WB___U154 ( .A(MEM_WB__n111), .Y(MEM_WB_ALU_result[7]) );
  BUFx3_ASAP7_75t_R MEM_WB___U155 ( .A(MEM_WB__n36), .Y(MEM_WB__n111) );
  BUFx2_ASAP7_75t_R MEM_WB___U156 ( .A(MEM_WB__n339), .Y(MEM_WB__n113) );
  BUFx3_ASAP7_75t_R MEM_WB___U157 ( .A(MEM_WB__n113), .Y(MEM_WB__n169) );
  BUFx2_ASAP7_75t_R MEM_WB___U158 ( .A(MEM_WB__n337), .Y(MEM_WB__n116) );
  BUFx2_ASAP7_75t_R MEM_WB___U159 ( .A(MEM_WB__n345), .Y(MEM_WB__n117) );
  BUFx3_ASAP7_75t_R MEM_WB___U160 ( .A(MEM_WB__n119), .Y(mem_data_out[21]) );
  BUFx2_ASAP7_75t_R MEM_WB___U161 ( .A(MEM_WB__n294), .Y(MEM_WB__n119) );
  BUFx2_ASAP7_75t_R MEM_WB___U162 ( .A(MEM_WB__n309), .Y(MEM_WB__n121) );
  BUFx2_ASAP7_75t_R MEM_WB___U163 ( .A(MEM_WB__n217), .Y(MEM_WB__n122) );
  INVx4_ASAP7_75t_R MEM_WB___U164 ( .A(MEM_mem_data[26]), .Y(MEM_WB__n258) );
  INVx4_ASAP7_75t_R MEM_WB___U165 ( .A(MEM_mem_data[24]), .Y(MEM_WB__n260) );
  BUFx2_ASAP7_75t_R MEM_WB___U166 ( .A(MEM_WB__n299), .Y(MEM_WB__n123) );
  BUFx2_ASAP7_75t_R MEM_WB___U167 ( .A(MEM_WB__n308), .Y(MEM_WB__n125) );
  BUFx2_ASAP7_75t_R MEM_WB___U168 ( .A(MEM_WB__n313), .Y(MEM_WB__n126) );
  BUFx3_ASAP7_75t_R MEM_WB___U169 ( .A(MEM_WB__n116), .Y(MEM_WB__n132) );
  BUFx4f_ASAP7_75t_R MEM_WB___U170 ( .A(MEM_WB__n136), .Y(mem_data_out[23]) );
  BUFx3_ASAP7_75t_R MEM_WB___U171 ( .A(MEM_WB__n39), .Y(MEM_WB__n136) );
  BUFx3_ASAP7_75t_R MEM_WB___U172 ( .A(MEM_WB__n40), .Y(MEM_WB__n138) );
  BUFx3_ASAP7_75t_R MEM_WB___U173 ( .A(MEM_WB__n27), .Y(MEM_WB__n140) );
  BUFx4f_ASAP7_75t_R MEM_WB___U174 ( .A(MEM_WB__n146), .Y(MEM_WB_ALU_result[30]) );
  BUFx3_ASAP7_75t_R MEM_WB___U175 ( .A(MEM_WB__n43), .Y(MEM_WB__n146) );
  BUFx4f_ASAP7_75t_R MEM_WB___U176 ( .A(MEM_WB__n148), .Y(MEM_WB_ALU_result[28]) );
  BUFx3_ASAP7_75t_R MEM_WB___U177 ( .A(MEM_WB__n8), .Y(MEM_WB__n148) );
  BUFx3_ASAP7_75t_R MEM_WB___U178 ( .A(MEM_WB__n102), .Y(MEM_WB__n150) );
  BUFx4f_ASAP7_75t_R MEM_WB___U179 ( .A(MEM_WB__n152), .Y(MEM_WB_ALU_result[14]) );
  BUFx3_ASAP7_75t_R MEM_WB___U180 ( .A(MEM_WB__n44), .Y(MEM_WB__n152) );
  BUFx4f_ASAP7_75t_R MEM_WB___U181 ( .A(MEM_WB__n154), .Y(MEM_WB_ALU_result[4]) );
  BUFx3_ASAP7_75t_R MEM_WB___U182 ( .A(MEM_WB__n104), .Y(MEM_WB__n154) );
  BUFx2_ASAP7_75t_R MEM_WB___U183 ( .A(MEM_WB__n214), .Y(MEM_WB__n155) );
  BUFx2_ASAP7_75t_R MEM_WB___U184 ( .A(MEM_WB__n215), .Y(MEM_WB__n156) );
  BUFx2_ASAP7_75t_R MEM_WB___U185 ( .A(MEM_WB__n213), .Y(MEM_WB__n157) );
  INVx4_ASAP7_75t_R MEM_WB___U186 ( .A(MEM_mem_data[31]), .Y(MEM_WB__n253) );
  INVx4_ASAP7_75t_R MEM_WB___U187 ( .A(MEM_mem_data[23]), .Y(MEM_WB__n261) );
  INVx4_ASAP7_75t_R MEM_WB___U188 ( .A(MEM_mem_data[22]), .Y(MEM_WB__n262) );
  INVx4_ASAP7_75t_R MEM_WB___U189 ( .A(MEM_mem_data[20]), .Y(MEM_WB__n264) );
  INVx4_ASAP7_75t_R MEM_WB___U190 ( .A(MEM_mem_data[18]), .Y(MEM_WB__n266) );
  INVx4_ASAP7_75t_R MEM_WB___U191 ( .A(MEM_mem_data[16]), .Y(MEM_WB__n268) );
  INVx4_ASAP7_75t_R MEM_WB___U192 ( .A(MEM_mem_data[15]), .Y(MEM_WB__n269) );
  INVx4_ASAP7_75t_R MEM_WB___U193 ( .A(MEM_mem_data[13]), .Y(MEM_WB__n271) );
  INVx4_ASAP7_75t_R MEM_WB___U194 ( .A(MEM_mem_data[9]), .Y(MEM_WB__n275) );
  INVx4_ASAP7_75t_R MEM_WB___U195 ( .A(MEM_mem_data[8]), .Y(MEM_WB__n276) );
  INVx4_ASAP7_75t_R MEM_WB___U196 ( .A(MEM_mem_data[6]), .Y(MEM_WB__n278) );
  INVx4_ASAP7_75t_R MEM_WB___U197 ( .A(MEM_mem_data[4]), .Y(MEM_WB__n280) );
  INVx4_ASAP7_75t_R MEM_WB___U198 ( .A(MEM_mem_data[2]), .Y(MEM_WB__n282) );
  INVx4_ASAP7_75t_R MEM_WB___U199 ( .A(MEM_mem_data[0]), .Y(MEM_WB__n284) );
  BUFx4f_ASAP7_75t_R MEM_WB___U200 ( .A(MEM_WB__n159), .Y(MEM_WB_ALU_result[22]) );
  BUFx3_ASAP7_75t_R MEM_WB___U201 ( .A(MEM_WB__n115), .Y(MEM_WB__n161) );
  BUFx3_ASAP7_75t_R MEM_WB___U202 ( .A(MEM_WB__n165), .Y(MEM_WB__n164) );
  BUFx2_ASAP7_75t_R MEM_WB___U203 ( .A(MEM_WB__n98), .Y(MEM_WB__n165) );
  BUFx3_ASAP7_75t_R MEM_WB___U204 ( .A(MEM_WB__n45), .Y(MEM_WB__n167) );
  BUFx4f_ASAP7_75t_R MEM_WB___U205 ( .A(MEM_WB__n171), .Y(mem_data_out[29]) );
  BUFx3_ASAP7_75t_R MEM_WB___U206 ( .A(MEM_WB__n15), .Y(MEM_WB__n171) );
  BUFx4f_ASAP7_75t_R MEM_WB___U207 ( .A(MEM_WB__n173), .Y(mem_data_out[26]) );
  BUFx3_ASAP7_75t_R MEM_WB___U208 ( .A(MEM_WB__n38), .Y(MEM_WB__n173) );
  BUFx4f_ASAP7_75t_R MEM_WB___U209 ( .A(MEM_WB__n175), .Y(mem_data_out[10]) );
  BUFx3_ASAP7_75t_R MEM_WB___U210 ( .A(MEM_WB__n6), .Y(MEM_WB__n175) );
  BUFx3_ASAP7_75t_R MEM_WB___U211 ( .A(MEM_WB__n47), .Y(MEM_WB__n177) );
  BUFx4f_ASAP7_75t_R MEM_WB___U212 ( .A(MEM_WB__n179), .Y(MEM_WB_ALU_result[2]) );
  BUFx3_ASAP7_75t_R MEM_WB___U213 ( .A(MEM_WB__n105), .Y(MEM_WB__n179) );
  BUFx4f_ASAP7_75t_R MEM_WB___U214 ( .A(MEM_WB__n183), .Y(MEM_WB_ALU_result[0]) );
  BUFx3_ASAP7_75t_R MEM_WB___U215 ( .A(MEM_WB__n117), .Y(MEM_WB__n183) );
  INVx4_ASAP7_75t_R MEM_WB___U216 ( .A(MEM_mem_data[30]), .Y(MEM_WB__n254) );
  INVx4_ASAP7_75t_R MEM_WB___U217 ( .A(MEM_mem_data[29]), .Y(MEM_WB__n255) );
  INVx4_ASAP7_75t_R MEM_WB___U218 ( .A(MEM_mem_data[28]), .Y(MEM_WB__n256) );
  INVx4_ASAP7_75t_R MEM_WB___U219 ( .A(MEM_mem_data[27]), .Y(MEM_WB__n257) );
  INVx4_ASAP7_75t_R MEM_WB___U220 ( .A(MEM_mem_data[25]), .Y(MEM_WB__n259) );
  INVx4_ASAP7_75t_R MEM_WB___U221 ( .A(MEM_mem_data[21]), .Y(MEM_WB__n263) );
  INVx4_ASAP7_75t_R MEM_WB___U222 ( .A(MEM_mem_data[19]), .Y(MEM_WB__n265) );
  INVx4_ASAP7_75t_R MEM_WB___U223 ( .A(MEM_mem_data[17]), .Y(MEM_WB__n267) );
  INVx4_ASAP7_75t_R MEM_WB___U224 ( .A(MEM_mem_data[14]), .Y(MEM_WB__n270) );
  INVx4_ASAP7_75t_R MEM_WB___U225 ( .A(MEM_mem_data[12]), .Y(MEM_WB__n272) );
  INVx4_ASAP7_75t_R MEM_WB___U226 ( .A(MEM_mem_data[11]), .Y(MEM_WB__n273) );
  INVx4_ASAP7_75t_R MEM_WB___U227 ( .A(MEM_mem_data[10]), .Y(MEM_WB__n274) );
  INVx4_ASAP7_75t_R MEM_WB___U228 ( .A(MEM_mem_data[7]), .Y(MEM_WB__n277) );
  INVx4_ASAP7_75t_R MEM_WB___U229 ( .A(MEM_mem_data[5]), .Y(MEM_WB__n279) );
  INVx4_ASAP7_75t_R MEM_WB___U230 ( .A(MEM_mem_data[3]), .Y(MEM_WB__n281) );
  INVx4_ASAP7_75t_R MEM_WB___U231 ( .A(MEM_mem_data[1]), .Y(MEM_WB__n283) );
  BUFx2_ASAP7_75t_R MEM_WB___U232 ( .A(EX_MEM_ALU_result[29]), .Y(MEM_WB__n221) );
  INVx1_ASAP7_75t_R MEM_WB___U233 ( .A(MEM_WB__n221), .Y(MEM_WB__n184) );
  BUFx2_ASAP7_75t_R MEM_WB___U234 ( .A(EX_MEM_ALU_result[25]), .Y(MEM_WB__n225) );
  INVx1_ASAP7_75t_R MEM_WB___U235 ( .A(MEM_WB__n225), .Y(MEM_WB__n185) );
  BUFx2_ASAP7_75t_R MEM_WB___U236 ( .A(EX_MEM_ALU_result[21]), .Y(MEM_WB__n229) );
  INVx1_ASAP7_75t_R MEM_WB___U237 ( .A(MEM_WB__n229), .Y(MEM_WB__n186) );
  BUFx2_ASAP7_75t_R MEM_WB___U238 ( .A(EX_MEM_ALU_result[17]), .Y(MEM_WB__n233) );
  INVx1_ASAP7_75t_R MEM_WB___U239 ( .A(MEM_WB__n233), .Y(MEM_WB__n187) );
  BUFx2_ASAP7_75t_R MEM_WB___U240 ( .A(EX_MEM_ALU_result[10]), .Y(MEM_WB__n240) );
  INVx1_ASAP7_75t_R MEM_WB___U241 ( .A(MEM_WB__n240), .Y(MEM_WB__n188) );
  BUFx2_ASAP7_75t_R MEM_WB___U242 ( .A(EX_MEM_ALU_result[5]), .Y(MEM_WB__n245) );
  INVx1_ASAP7_75t_R MEM_WB___U243 ( .A(MEM_WB__n245), .Y(MEM_WB__n189) );
  BUFx3_ASAP7_75t_R MEM_WB___U244 ( .A(MEM_WB__n197), .Y(mem_data_out[15]) );
  BUFx2_ASAP7_75t_R MEM_WB___U245 ( .A(MEM_WB__n123), .Y(MEM_WB__n197) );
  BUFx3_ASAP7_75t_R MEM_WB___U246 ( .A(MEM_WB__n203), .Y(mem_data_out[6]) );
  BUFx2_ASAP7_75t_R MEM_WB___U247 ( .A(MEM_WB__n125), .Y(MEM_WB__n203) );
  BUFx4f_ASAP7_75t_R MEM_WB___U248 ( .A(MEM_WB__n205), .Y(mem_data_out[31]) );
  BUFx3_ASAP7_75t_R MEM_WB___U249 ( .A(MEM_WB__n13), .Y(MEM_WB__n205) );
  BUFx3_ASAP7_75t_R MEM_WB___U250 ( .A(MEM_WB__n19), .Y(MEM_WB__n207) );
  BUFx3_ASAP7_75t_R MEM_WB___U251 ( .A(MEM_WB__n114), .Y(MEM_WB__n209) );
  INVx1_ASAP7_75t_R MEM_WB___U252 ( .A(MEM_WB__n64), .Y(MEM_WB__n217) );
  INVx1_ASAP7_75t_R MEM_WB___U253 ( .A(EX_MEM_rd[1]), .Y(MEM_WB__n216) );
  INVx1_ASAP7_75t_R MEM_WB___U254 ( .A(MEM_WB__n107), .Y(MEM_WB__n215) );
  INVx1_ASAP7_75t_R MEM_WB___U255 ( .A(MEM_WB__n49), .Y(MEM_WB__n214) );
  INVx1_ASAP7_75t_R MEM_WB___U256 ( .A(MEM_WB__n106), .Y(MEM_WB__n213) );
  INVx1_ASAP7_75t_R MEM_WB___U257 ( .A(EX_MEM_ALU_result[0]), .Y(MEM_WB__n250) );
  INVx1_ASAP7_75t_R MEM_WB___U258 ( .A(EX_MEM_ALU_result[1]), .Y(MEM_WB__n249) );
  INVx1_ASAP7_75t_R MEM_WB___U259 ( .A(EX_MEM_ALU_result[2]), .Y(MEM_WB__n248) );
  INVx1_ASAP7_75t_R MEM_WB___U260 ( .A(EX_MEM_ALU_result[3]), .Y(MEM_WB__n247) );
  INVx1_ASAP7_75t_R MEM_WB___U261 ( .A(EX_MEM_ALU_result[4]), .Y(MEM_WB__n246) );
  INVx1_ASAP7_75t_R MEM_WB___U262 ( .A(EX_MEM_ALU_result[6]), .Y(MEM_WB__n244) );
  INVx1_ASAP7_75t_R MEM_WB___U263 ( .A(EX_MEM_ALU_result[7]), .Y(MEM_WB__n243) );
  INVx1_ASAP7_75t_R MEM_WB___U264 ( .A(EX_MEM_ALU_result[8]), .Y(MEM_WB__n242) );
  INVx1_ASAP7_75t_R MEM_WB___U265 ( .A(EX_MEM_ALU_result[9]), .Y(MEM_WB__n241) );
  INVx1_ASAP7_75t_R MEM_WB___U266 ( .A(EX_MEM_ALU_result[11]), .Y(MEM_WB__n239) );
  INVx1_ASAP7_75t_R MEM_WB___U267 ( .A(EX_MEM_ALU_result[12]), .Y(MEM_WB__n238) );
  INVx1_ASAP7_75t_R MEM_WB___U268 ( .A(EX_MEM_ALU_result[13]), .Y(MEM_WB__n237) );
  INVx1_ASAP7_75t_R MEM_WB___U269 ( .A(EX_MEM_ALU_result[14]), .Y(MEM_WB__n236) );
  INVx1_ASAP7_75t_R MEM_WB___U270 ( .A(EX_MEM_ALU_result[15]), .Y(MEM_WB__n235) );
  INVx1_ASAP7_75t_R MEM_WB___U271 ( .A(EX_MEM_ALU_result[16]), .Y(MEM_WB__n234) );
  INVx1_ASAP7_75t_R MEM_WB___U272 ( .A(EX_MEM_ALU_result[18]), .Y(MEM_WB__n232) );
  INVx1_ASAP7_75t_R MEM_WB___U273 ( .A(EX_MEM_ALU_result[19]), .Y(MEM_WB__n231) );
  INVx1_ASAP7_75t_R MEM_WB___U274 ( .A(EX_MEM_ALU_result[20]), .Y(MEM_WB__n230) );
  INVx1_ASAP7_75t_R MEM_WB___U275 ( .A(EX_MEM_ALU_result[22]), .Y(MEM_WB__n228) );
  INVx1_ASAP7_75t_R MEM_WB___U276 ( .A(EX_MEM_ALU_result[23]), .Y(MEM_WB__n227) );
  INVx1_ASAP7_75t_R MEM_WB___U277 ( .A(EX_MEM_ALU_result[24]), .Y(MEM_WB__n226) );
  INVx1_ASAP7_75t_R MEM_WB___U278 ( .A(EX_MEM_ALU_result[26]), .Y(MEM_WB__n224) );
  INVx1_ASAP7_75t_R MEM_WB___U279 ( .A(EX_MEM_ALU_result[27]), .Y(MEM_WB__n223) );
  INVx1_ASAP7_75t_R MEM_WB___U280 ( .A(EX_MEM_ALU_result[28]), .Y(MEM_WB__n222) );
  INVx1_ASAP7_75t_R MEM_WB___U281 ( .A(EX_MEM_ALU_result[30]), .Y(MEM_WB__n220) );
  INVx1_ASAP7_75t_R MEM_WB___U282 ( .A(EX_MEM_ALU_result[31]), .Y(MEM_WB__n219) );
  INVx1_ASAP7_75t_R MEM_WB___U283 ( .A(EX_MEM_MemRead), .Y(MEM_WB__n251) );
  INVx1_ASAP7_75t_R MEM_WB___U284 ( .A(EX_MEM_MemToReg), .Y(MEM_WB__n252) );
  INVx1_ASAP7_75t_R MEM_WB___U285 ( .A(EX_MEM_RegWrite), .Y(MEM_WB__n218) );

    OA22x2_ASAP7_75t_R WB___U1 ( .A1(WB__n11), .A2(WB__n88), .B1(WB__n12), .B2(WB__n56), .Y(WB__n101) );
  INVx2_ASAP7_75t_R WB___U2 ( .A(WB__n101), .Y(WB_write_back_data[0]) );
  BUFx4f_ASAP7_75t_R WB___U3 ( .A(MEM_WB_rd[1]), .Y(WB_rd[1]) );
  BUFx3_ASAP7_75t_R WB___U4 ( .A(WB__n47), .Y(WB__n61) );
  INVx1_ASAP7_75t_R WB___U5 ( .A(WB__n47), .Y(WB__n85) );
  INVx1_ASAP7_75t_R WB___U6 ( .A(WB__n47), .Y(WB__n94) );
  INVx1_ASAP7_75t_R WB___U7 ( .A(WB__n83), .Y(WB__n76) );
  INVxp67_ASAP7_75t_R WB___U8 ( .A(WB__n3), .Y(WB__n2) );
  INVxp33_ASAP7_75t_R WB___U9 ( .A(WB__n95), .Y(WB__n26) );
  INVx2_ASAP7_75t_R WB___U10 ( .A(WB__n48), .Y(WB__n47) );
  INVx1_ASAP7_75t_R WB___U11 ( .A(WB__n57), .Y(WB__n48) );
  AO22x2_ASAP7_75t_R WB___U12 ( .A1(MEM_WB_ALU_result[31]), .A2(WB__n3), .B1(MEM_WB_mem_data[31]), 
        .B2(WB__n94), .Y(WB_write_back_data[31]) );
  BUFx2_ASAP7_75t_R WB___U13 ( .A(WB__n47), .Y(WB__n3) );
  NAND2xp5_ASAP7_75t_R WB___U14 ( .A(MEM_WB_mem_data[8]), .B(WB__n89), .Y(WB__n54) );
  INVx1_ASAP7_75t_R WB___U15 ( .A(WB__n83), .Y(WB__n75) );
  AO22x2_ASAP7_75t_R WB___U16 ( .A1(MEM_WB_ALU_result[26]), .A2(WB__n63), .B1(MEM_WB_mem_data[26]), 
        .B2(WB__n86), .Y(WB_write_back_data[26]) );
  INVx1_ASAP7_75t_R WB___U17 ( .A(WB__n83), .Y(WB__n77) );
  INVxp33_ASAP7_75t_R WB___U18 ( .A(MEM_WB_ALU_result[2]), .Y(WB__n18) );
  INVxp67_ASAP7_75t_R WB___U19 ( .A(WB__n96), .Y(WB__n17) );
  INVxp67_ASAP7_75t_R WB___U20 ( .A(WB__n96), .Y(WB__n87) );
  NOR2xp67_ASAP7_75t_R WB___U21 ( .A(WB__n35), .B(WB__n80), .Y(WB__n14) );
  INVx2_ASAP7_75t_R WB___U22 ( .A(WB__n95), .Y(WB__n88) );
  OAI22xp33_ASAP7_75t_R WB___U23 ( .A1(WB__n39), .A2(WB__n87), .B1(WB__n40), .B2(WB__n67), .Y(
        WB_write_back_data[13]) );
  BUFx2_ASAP7_75t_R WB___U24 ( .A(WB__n58), .Y(WB__n95) );
  NAND2xp33_ASAP7_75t_R WB___U25 ( .A(MEM_WB_ALU_result[9]), .B(WB__n76), .Y(WB__n4) );
  NAND2xp5_ASAP7_75t_R WB___U26 ( .A(MEM_WB_mem_data[9]), .B(WB__n38), .Y(WB__n5) );
  NAND2xp67_ASAP7_75t_R WB___U27 ( .A(WB__n4), .B(WB__n5), .Y(WB_write_back_data[9]) );
  OAI22xp33_ASAP7_75t_R WB___U28 ( .A1(WB__n17), .A2(WB__n31), .B1(WB__n32), .B2(WB__n66), .Y(
        WB_write_back_data[22]) );
  OAI22xp5_ASAP7_75t_R WB___U29 ( .A1(WB__n15), .A2(WB__n89), .B1(WB__n16), .B2(WB__n66), .Y(
        WB_write_back_data[27]) );
  AO22x1_ASAP7_75t_R WB___U30 ( .A1(MEM_WB_ALU_result[20]), .A2(WB__n95), .B1(MEM_WB_mem_data[20]), 
        .B2(WB__n94), .Y(WB_write_back_data[20]) );
  HB1xp67_ASAP7_75t_R WB___U31 ( .A(WB__n96), .Y(WB__n66) );
  INVxp33_ASAP7_75t_R WB___U32 ( .A(WB__n96), .Y(WB__n90) );
  OAI22xp5_ASAP7_75t_R WB___U33 ( .A1(WB__n43), .A2(WB__n87), .B1(WB__n44), .B2(WB__n81), .Y(
        WB_write_back_data[25]) );
  INVx5_ASAP7_75t_R WB___U34 ( .A(WB__n56), .Y(WB__n89) );
  INVxp67_ASAP7_75t_R WB___U35 ( .A(MEM_WB_mem_data[13]), .Y(WB__n40) );
  INVx1_ASAP7_75t_R WB___U36 ( .A(WB__n87), .Y(WB__n78) );
  INVxp33_ASAP7_75t_R WB___U37 ( .A(WB__n96), .Y(WB__n84) );
  NOR2xp67_ASAP7_75t_R WB___U38 ( .A(WB__n34), .B(WB__n17), .Y(WB__n13) );
  INVx1_ASAP7_75t_R WB___U39 ( .A(WB__n67), .Y(WB__n86) );
  BUFx2_ASAP7_75t_R WB___U40 ( .A(WB__n58), .Y(WB__n67) );
  INVx1_ASAP7_75t_R WB___U41 ( .A(MEM_WB_ALU_result[0]), .Y(WB__n11) );
  INVx1_ASAP7_75t_R WB___U42 ( .A(MEM_WB_ALU_result[13]), .Y(WB__n39) );
  OAI22xp33_ASAP7_75t_R WB___U43 ( .A1(WB__n83), .A2(WB__n18), .B1(WB__n19), .B2(WB__n56), .Y(
        WB_write_back_data[2]) );
  NAND2xp67_ASAP7_75t_R WB___U44 ( .A(WB__n20), .B(WB__n21), .Y(WB_write_back_data[1]) );
  INVx2_ASAP7_75t_R WB___U45 ( .A(WB__n88), .Y(WB__n81) );
  OAI22xp5_ASAP7_75t_R WB___U46 ( .A1(WB__n41), .A2(WB__n89), .B1(WB__n42), .B2(WB__n78), .Y(WB__n99)
         );
  INVxp33_ASAP7_75t_R WB___U47 ( .A(MEM_WB_ALU_result[24]), .Y(WB__n9) );
  OAI22xp33_ASAP7_75t_R WB___U48 ( .A1(WB__n51), .A2(WB__n90), .B1(WB__n52), .B2(WB__n3), .Y(
        WB_write_back_data[17]) );
  NAND2x1_ASAP7_75t_R WB___U49 ( .A(WB__n36), .B(WB__n37), .Y(WB_write_back_data[21]) );
  NAND2xp5_ASAP7_75t_R WB___U50 ( .A(MEM_WB_mem_data[1]), .B(WB__n85), .Y(WB__n21) );
  INVx1_ASAP7_75t_R WB___U51 ( .A(WB__n89), .Y(WB__n63) );
  NAND2xp33_ASAP7_75t_R WB___U52 ( .A(MEM_WB_ALU_result[3]), .B(WB__n67), .Y(WB__n7) );
  NAND2xp33_ASAP7_75t_R WB___U53 ( .A(MEM_WB_mem_data[3]), .B(WB__WB__n86), .Y(WB__n8) );
  NAND2xp67_ASAP7_75t_R WB___U54 ( .A(WB__n7), .B(WB__n8), .Y(WB_write_back_data[3]) );
  NAND2xp5_ASAP7_75t_R WB___U55 ( .A(MEM_WB_ALU_result[1]), .B(WB__n96), .Y(WB__n20) );
  NOR2xp33_ASAP7_75t_R WB___U56 ( .A(WB__n30), .B(WB__n76), .Y(WB__n25) );
  INVxp67_ASAP7_75t_R WB___U57 ( .A(MEM_WB_mem_data[24]), .Y(WB__n10) );
  OAI22xp33_ASAP7_75t_R WB___U58 ( .A1(WB__n9), .A2(WB__n2), .B1(WB__n10), .B2(WB__n75), .Y(
        WB_write_back_data[24]) );
  NAND2xp5_ASAP7_75t_R WB___U59 ( .A(MEM_WB_mem_data[6]), .B(WB__n86), .Y(WB__n23) );
  INVxp67_ASAP7_75t_R WB___U60 ( .A(WB__n67), .Y(WB__n93) );
  OAI22xp33_ASAP7_75t_R WB___U61 ( .A1(WB__n49), .A2(WB__n93), .B1(WB__n50), .B2(WB__n67), .Y(
        WB_write_back_data[14]) );
  NAND2x1p5_ASAP7_75t_R WB___U62 ( .A(MEM_WB_ALU_result[21]), .B(WB__n81), .Y(WB__n36) );
  BUFx3_ASAP7_75t_R WB___U63 ( .A(WB__n99), .Y(WB_write_back_data[5]) );
  INVx2_ASAP7_75t_R WB___U64 ( .A(WB__n64), .Y(WB_write_back_data[11]) );
  BUFx6f_ASAP7_75t_R WB___U65 ( .A(WB__n100), .Y(WB_write_back_data[4]) );
  CKINVDCx20_ASAP7_75t_R WB___U66 ( .A(MEM_WB_mem_data[0]), .Y(WB__n12) );
  NAND2xp33_ASAP7_75t_R WB___U67 ( .A(MEM_WB_ALU_result[8]), .B(WB__n56), .Y(WB__n53) );
  OR2x2_ASAP7_75t_R WB___U68 ( .A(WB__n13), .B(WB__n14), .Y(WB_write_back_data[19]) );
  INVx1_ASAP7_75t_R WB___U69 ( .A(MEM_WB_ALU_result[19]), .Y(WB__n34) );
  INVxp67_ASAP7_75t_R WB___U70 ( .A(MEM_WB_mem_data[19]), .Y(WB__n35) );
  INVx1_ASAP7_75t_R WB___U71 ( .A(WB__n85), .Y(WB__n80) );
  BUFx4f_ASAP7_75t_R WB___U72 ( .A(WB__n98), .Y(WB_write_back_data[12]) );
  INVx2_ASAP7_75t_R WB___U73 ( .A(MEM_WB_mem_data[2]), .Y(WB__n19) );
  CKINVDCx20_ASAP7_75t_R WB___U74 ( .A(MEM_WB_ALU_result[27]), .Y(WB__n15) );
  CKINVDCx20_ASAP7_75t_R WB___U75 ( .A(MEM_WB_mem_data[27]), .Y(WB__n16) );
  BUFx2_ASAP7_75t_R WB___U76 ( .A(WB__n33), .Y(WB__n64) );
  BUFx12f_ASAP7_75t_R WB___U77 ( .A(n51), .Y(WB_rd[2]) );
  INVx1_ASAP7_75t_R WB___U78 ( .A(MEM_WB_mem_data[23]), .Y(WB__n28) );
  NAND2xp33_ASAP7_75t_R WB___U79 ( .A(WB__n53), .B(WB__n54), .Y(WB_write_back_data[8]) );
  NAND2xp67_ASAP7_75t_R WB___U80 ( .A(WB__n22), .B(WB__n23), .Y(WB_write_back_data[6]) );
  AOI22xp33_ASAP7_75t_R WB___U81 ( .A1(MEM_WB_ALU_result[11]), .A2(WB__n80), .B1(MEM_WB_mem_data[11]), 
        .B2(WB__n17), .Y(WB__n33) );
  BUFx3_ASAP7_75t_R WB___U82 ( .A(WB__n82), .Y(WB__n83) );
  INVxp33_ASAP7_75t_R WB___U83 ( .A(MEM_WB_ALU_result[22]), .Y(WB__n31) );
  INVx1_ASAP7_75t_R WB___U84 ( .A(MEM_WB_ALU_result[5]), .Y(WB__n41) );
  INVx1_ASAP7_75t_R WB___U85 ( .A(WB__n89), .Y(WB__n79) );
  INVxp33_ASAP7_75t_R WB___U86 ( .A(WB__n80), .Y(WB__n38) );
  BUFx3_ASAP7_75t_R WB___U87 ( .A(MEM_WB_rd[4]), .Y(WB_rd[4]) );
  HB1xp67_ASAP7_75t_R WB___U88 ( .A(WB__n97), .Y(WB_write_back_data[23]) );
  INVxp67_ASAP7_75t_R WB___U89 ( .A(MEM_WB_ALU_result[23]), .Y(WB__n27) );
  INVxp67_ASAP7_75t_R WB___U90 ( .A(WB__n79), .Y(WB__n92) );
  BUFx3_ASAP7_75t_R WB___U91 ( .A(MEM_WB_rd[3]), .Y(WB_rd[3]) );
  NAND2xp33_ASAP7_75t_R WB___U92 ( .A(MEM_WB_mem_data[21]), .B(WB__n2), .Y(WB__n37) );
  AO22x1_ASAP7_75t_R WB___U93 ( .A1(MEM_WB_ALU_result[30]), .A2(WB__n3), .B1(MEM_WB_mem_data[30]), 
        .B2(WB__n94), .Y(WB_write_back_data[30]) );
  BUFx6f_ASAP7_75t_R WB___U94 ( .A(WB__n61), .Y(WB__n56) );
  INVxp67_ASAP7_75t_R WB___U95 ( .A(MEM_WB_mem_data[5]), .Y(WB__n42) );
  AO22x1_ASAP7_75t_R WB___U96 ( .A1(MEM_WB_ALU_result[15]), .A2(WB__n79), .B1(MEM_WB_mem_data[15]), 
        .B2(WB__n91), .Y(WB_write_back_data[15]) );
  INVxp67_ASAP7_75t_R WB___U97 ( .A(WB__n62), .Y(WB__n91) );
  NAND2xp5_ASAP7_75t_R WB___U98 ( .A(MEM_WB_ALU_result[6]), .B(WB__n78), .Y(WB__n22) );
  NOR2xp33_ASAP7_75t_R WB___U99 ( .A(WB__n29), .B(WB__n94), .Y(WB__n24) );
  OR2x2_ASAP7_75t_R WB___U100 ( .A(WB__n24), .B(WB__n25), .Y(WB__n100) );
  INVxp33_ASAP7_75t_R WB___U101 ( .A(MEM_WB_ALU_result[4]), .Y(WB__n29) );
  INVxp33_ASAP7_75t_R WB___U102 ( .A(MEM_WB_mem_data[4]), .Y(WB__n30) );
  INVxp33_ASAP7_75t_R WB___U103 ( .A(MEM_WB_mem_data[22]), .Y(WB__n32) );
  OAI22xp33_ASAP7_75t_R WB___U104 ( .A1(WB__n27), .A2(WB__n83), .B1(WB__n28), .B2(WB__n67), .Y(WB__n97)
         );
  OAI22xp33_ASAP7_75t_R WB___U105 ( .A1(WB__n45), .A2(WB__n83), .B1(WB__n46), .B2(WB__n81), .Y(
        WB_write_back_data[29]) );
  BUFx12f_ASAP7_75t_R WB___U106 ( .A(MEM_WB_rd[0]), .Y(WB_rd[0]) );
  INVx2_ASAP7_75t_R WB___U107 ( .A(MEM_WB_mem_data[17]), .Y(WB__n52) );
  INVx1_ASAP7_75t_R WB___U108 ( .A(n14), .Y(WB__n44) );
  AO22x1_ASAP7_75t_R WB___U109 ( .A1(MEM_WB_ALU_result[12]), .A2(WB__n75), .B1(MEM_WB_mem_data[12]), 
        .B2(WB__n84), .Y(WB__n98) );
  CKINVDCx20_ASAP7_75t_R WB___U110 ( .A(MEM_WB_ALU_result[25]), .Y(WB__n43) );
  HB1xp67_ASAP7_75t_R WB___U111 ( .A(WB__n78), .Y(WB__n62) );
  HB1xp67_ASAP7_75t_R WB___U112 ( .A(WB__n26), .Y(WB__n55) );
  CKINVDCx20_ASAP7_75t_R WB___U113 ( .A(MEM_WB_ALU_result[29]), .Y(WB__n45) );
  CKINVDCx20_ASAP7_75t_R WB___U114 ( .A(MEM_WB_mem_data[29]), .Y(WB__n46) );
  HB1xp67_ASAP7_75t_R WB___U115 ( .A(WB__n48), .Y(WB__n82) );
  HB1xp67_ASAP7_75t_R WB___U116 ( .A(WB__n57), .Y(WB__n58) );
  INVx1_ASAP7_75t_R WB___U117 ( .A(MEM_WB_MemtoReg), .Y(WB__n57) );
  AO22x1_ASAP7_75t_R WB___U118 ( .A1(MEM_WB_ALU_result[28]), .A2(WB__n80), .B1(MEM_WB_mem_data[28]), 
        .B2(WB__n55), .Y(WB_write_back_data[28]) );
  INVx1_ASAP7_75t_R WB___U119 ( .A(MEM_WB_mem_data[14]), .Y(WB__n50) );
  INVx1_ASAP7_75t_R WB___U120 ( .A(MEM_WB_ALU_result[17]), .Y(WB__n51) );
  INVx1_ASAP7_75t_R WB___U121 ( .A(MEM_WB_ALU_result[14]), .Y(WB__n49) );
  HB1xp67_ASAP7_75t_R WB___U122 ( .A(WB__n57), .Y(WB__n96) );
  AO22x1_ASAP7_75t_R WB___U123 ( .A1(MEM_WB_ALU_result[10]), .A2(WB__n77), .B1(MEM_WB_mem_data[10]), 
        .B2(WB__n84), .Y(WB_write_back_data[10]) );
  AO22x1_ASAP7_75t_R WB___U124 ( .A1(MEM_WB_ALU_result[7]), .A2(WB__n67), .B1(MEM_WB_mem_data[7]), 
        .B2(WB__n88), .Y(WB_write_back_data[7]) );
  AO22x1_ASAP7_75t_R WB___U125 ( .A1(MEM_WB_ALU_result[18]), .A2(WB__n80), .B1(MEM_WB_mem_data[18]), 
        .B2(WB__n17), .Y(WB_write_back_data[18]) );
  AO22x1_ASAP7_75t_R WB___U126 ( .A1(MEM_WB_ALU_result[16]), .A2(WB__n80), .B1(MEM_WB_mem_data[16]), 
        .B2(WB__n92), .Y(WB_write_back_data[16]) );
 
  DHLx3_ASAP7_75t_R FORWARDING___ForwardA_reg_0_ ( .CLK(FORWARDING__n118), .D(FORWARDING__n131), .Q(FORWARDING__n505) );
  DHLx3_ASAP7_75t_R FORWARDING___ForwardA_reg_1_ ( .CLK(FORWARDING__n118), .D(FORWARDING__n166), .Q(FORWARDING__n504) );
  DHLx3_ASAP7_75t_R FORWARDING___ForwardB_reg_1_ ( .CLK(FORWARDING__n118), .D(FORWARDING__n63), .Q(FORWARDING__n506) );
  DHLx3_ASAP7_75t_R FORWARDING___ForwardB_reg_0_ ( .CLK(FORWARDING__n118), .D(FORWARDING__n122), .Q(FORWARDING__n507) );
  CKINVDCx5p33_ASAP7_75t_R FORWARDING___U3 ( .A(FORWARDING__n361), .Y(FORWARDING__n23) );
  CKINVDCx20_ASAP7_75t_R FORWARDING___U4 ( .A(FORWARDING__n406), .Y(FORWARDING__n244) );
  BUFx16f_ASAP7_75t_R FORWARDING___U5 ( .A(MEM_WB_ALU_result[15]), .Y(FORWARDING__n406) );
  INVx4_ASAP7_75t_R FORWARDING___U6 ( .A(FORWARDING__n270), .Y(forwarding_MEM_WB[26]) );
  BUFx6f_ASAP7_75t_R FORWARDING___U7 ( .A(FORWARDING__n316), .Y(FORWARDING__n270) );
  BUFx4f_ASAP7_75t_R FORWARDING___U8 ( .A(FORWARDING__n374), .Y(FORWARDING__n72) );
  HB1xp67_ASAP7_75t_R FORWARDING___U9 ( .A(FORWARDING__n36), .Y(FORWARDING__FORWARDING__n369) );
  BUFx2_ASAP7_75t_R FORWARDING___U10 ( .A(FORWARDING__n37), .Y(FORWARDING__n73) );
  BUFx4f_ASAP7_75t_R FORWARDING___U11 ( .A(FORWARDING__n37), .Y(FORWARDING__n40) );
  BUFx6f_ASAP7_75t_R FORWARDING___U12 ( .A(FORWARDING__n360), .Y(FORWARDING__n97) );
  BUFx4f_ASAP7_75t_R FORWARDING___U13 ( .A(FORWARDING__n374), .Y(FORWARDING__n360) );
  AND2x4_ASAP7_75t_R FORWARDING___U14 ( .A(FORWARDING__n298), .B(FORWARDING__n365), .Y(FORWARDING__n401) );
  INVxp33_ASAP7_75t_R FORWARDING___U15 ( .A(FORWARDING__n139), .Y(forwarding_MEM_WB[1]) );
  BUFx3_ASAP7_75t_R FORWARDING___U16 ( .A(FORWARDING__n38), .Y(FORWARDING__n129) );
  INVx2_ASAP7_75t_R FORWARDING___U17 ( .A(MEM_WB_ALU_result[13]), .Y(FORWARDING__n402) );
  BUFx6f_ASAP7_75t_R FORWARDING___U18 ( .A(FORWARDING__n73), .Y(FORWARDING__n361) );
  HB1xp67_ASAP7_75t_R FORWARDING___U19 ( .A(FORWARDING__n37), .Y(FORWARDING__n36) );
  OAI21xp33_ASAP7_75t_R FORWARDING___U20 ( .A1(FORWARDING__n372), .A2(FORWARDING__n301), .B(FORWARDING__n76), .Y(
        forwarding_MEM_WB[20]) );
  INVxp33_ASAP7_75t_R FORWARDING___U21 ( .A(FORWARDING__n209), .Y(forwarding_MEM_WB[23]) );
  BUFx2_ASAP7_75t_R FORWARDING___U22 ( .A(FORWARDING__n36), .Y(FORWARDING__n39) );
  AND2x2_ASAP7_75t_R FORWARDING___U23 ( .A(MEM_WB_mem_data[23]), .B(FORWARDING__n369), .Y(FORWARDING__n421) );
  INVxp33_ASAP7_75t_R FORWARDING___U24 ( .A(FORWARDING__n362), .Y(FORWARDING__n17) );
  INVxp67_ASAP7_75t_R FORWARDING___U25 ( .A(MEM_WB_ALU_result[1]), .Y(FORWARDING__n379) );
  AND2x2_ASAP7_75t_R FORWARDING___U26 ( .A(MEM_WB_mem_data[1]), .B(FORWARDING__n129), .Y(FORWARDING__n378)
         );
  BUFx6f_ASAP7_75t_R FORWARDING___U27 ( .A(FORWARDING__n361), .Y(FORWARDING__n375) );
  HB1xp67_ASAP7_75t_R FORWARDING___U28 ( .A(FORWARDING__n72), .Y(FORWARDING__n363) );
  BUFx6f_ASAP7_75t_R FORWARDING___U29 ( .A(FORWARDING__n96), .Y(FORWARDING__n365) );
  INVx1_ASAP7_75t_R FORWARDING___U30 ( .A(FORWARDING__n365), .Y(FORWARDING__n12) );
  INVxp67_ASAP7_75t_R FORWARDING___U31 ( .A(FORWARDING__n224), .Y(forwarding_MEM_WB[22]) );
  AND2x2_ASAP7_75t_R FORWARDING___U32 ( .A(MEM_WB_mem_data[29]), .B(FORWARDING__n373), .Y(FORWARDING__n432) );
  HB1xp67_ASAP7_75t_R FORWARDING___U33 ( .A(FORWARDING__n373), .Y(FORWARDING__n366) );
  INVxp67_ASAP7_75t_R FORWARDING___U34 ( .A(FORWARDING__n476), .Y(FORWARDING__n2) );
  INVx1_ASAP7_75t_R FORWARDING___U35 ( .A(FORWARDING__n434), .Y(FORWARDING__n3) );
  AND2x2_ASAP7_75t_R FORWARDING___U36 ( .A(MEM_WB_mem_data[30]), .B(FORWARDING__n130), .Y(FORWARDING__n434) );
  BUFx6f_ASAP7_75t_R FORWARDING___U37 ( .A(FORWARDING__n39), .Y(FORWARDING__n130) );
  HB1xp67_ASAP7_75t_R FORWARDING___U38 ( .A(FORWARDING__n374), .Y(FORWARDING__n38) );
  BUFx3_ASAP7_75t_R FORWARDING___U39 ( .A(FORWARDING__n96), .Y(FORWARDING__n364) );
  BUFx4f_ASAP7_75t_R FORWARDING___U40 ( .A(FORWARDING__n97), .Y(FORWARDING__n96) );
  INVx4_ASAP7_75t_R FORWARDING___U41 ( .A(FORWARDING__n103), .Y(forwarding_MEM_WB[27]) );
  BUFx6f_ASAP7_75t_R FORWARDING___U42 ( .A(FORWARDING__n281), .Y(FORWARDING__n103) );
  INVx1_ASAP7_75t_R FORWARDING___U43 ( .A(FORWARDING__n81), .Y(forwarding_MEM_WB[11]) );
  BUFx6f_ASAP7_75t_R FORWARDING___U44 ( .A(FORWARDING__n40), .Y(FORWARDING__n373) );
  INVxp33_ASAP7_75t_R FORWARDING___U45 ( .A(FORWARDING__n202), .Y(forwarding_MEM_WB[3]) );
  BUFx2_ASAP7_75t_R FORWARDING___U46 ( .A(MEM_WB_MemRead), .Y(FORWARDING__n374) );
  BUFx2_ASAP7_75t_R FORWARDING___U47 ( .A(MEM_WB_MemRead), .Y(FORWARDING__n37) );
  BUFx3_ASAP7_75t_R FORWARDING___U48 ( .A(FORWARDING__n159), .Y(forwarding_MEM_WB[16]) );
  INVxp33_ASAP7_75t_R FORWARDING___U49 ( .A(FORWARDING__n150), .Y(FORWARDING__n308) );
  HB1xp67_ASAP7_75t_R FORWARDING___U50 ( .A(FORWARDING__n482), .Y(FORWARDING__n150) );
  HB1xp67_ASAP7_75t_R FORWARDING___U51 ( .A(FORWARDING__n308), .Y(forwarding_MEM_WB[24]) );
  INVxp67_ASAP7_75t_R FORWARDING___U52 ( .A(FORWARDING__n164), .Y(FORWARDING__n87) );
  HB1xp67_ASAP7_75t_R FORWARDING___U53 ( .A(FORWARDING__n425), .Y(FORWARDING__n164) );
  BUFx6f_ASAP7_75t_R FORWARDING___U54 ( .A(FORWARDING__n72), .Y(FORWARDING__n370) );
  INVx1_ASAP7_75t_R FORWARDING___U55 ( .A(FORWARDING__n475), .Y(forwarding_MEM_WB[31]) );
  NAND2xp33_ASAP7_75t_R FORWARDING___U56 ( .A(MEM_WB_mem_data[28]), .B(FORWARDING__n373), .Y(
        n5) );
  INVx2_ASAP7_75t_R FORWARDING___U57 ( .A(FORWARDING__n153), .Y(FORWARDING__n310) );
  INVx4_ASAP7_75t_R FORWARDING___U58 ( .A(FORWARDING__n61), .Y(forwarding_MEM_WB[25]) );
  BUFx12f_ASAP7_75t_R FORWARDING___U59 ( .A(FORWARDING__n130), .Y(FORWARDING__n358) );
  OAI21xp33_ASAP7_75t_R FORWARDING___U60 ( .A1(FORWARDING__n274), .A2(FORWARDING__n359), .B(FORWARDING__n98), .Y(
        forwarding_MEM_WB[19]) );
  INVx1_ASAP7_75t_R FORWARDING___U61 ( .A(FORWARDING__n110), .Y(forwarding_MEM_WB[6]) );
  HB1xp67_ASAP7_75t_R FORWARDING___U62 ( .A(MEM_WB_RegWrite), .Y(FORWARDING__n120) );
  INVx4_ASAP7_75t_R FORWARDING___U63 ( .A(MEM_WB_mem_data[5]), .Y(FORWARDING__n19) );
  INVx1_ASAP7_75t_R FORWARDING___U64 ( .A(FORWARDING__n386), .Y(FORWARDING__n6) );
  NOR2x1p5_ASAP7_75t_R FORWARDING___U65 ( .A(FORWARDING__n19), .B(FORWARDING__n23), .Y(FORWARDING__n386) );
  BUFx2_ASAP7_75t_R FORWARDING___U66 ( .A(FORWARDING__n72), .Y(FORWARDING__n362) );
  BUFx6f_ASAP7_75t_R FORWARDING___U67 ( .A(FORWARDING__n129), .Y(FORWARDING__n359) );
  HB1xp67_ASAP7_75t_R FORWARDING___U68 ( .A(FORWARDING__n210), .Y(FORWARDING__n209) );
  INVxp67_ASAP7_75t_R FORWARDING___U69 ( .A(FORWARDING__n22), .Y(FORWARDING__n489) );
  HB1xp67_ASAP7_75t_R FORWARDING___U70 ( .A(FORWARDING__n483), .Y(FORWARDING__n210) );
  INVx2_ASAP7_75t_R FORWARDING___U71 ( .A(FORWARDING__n421), .Y(FORWARDING__n320) );
  INVxp33_ASAP7_75t_R FORWARDING___U72 ( .A(FORWARDING__n264), .Y(FORWARDING__n201) );
  HB1xp67_ASAP7_75t_R FORWARDING___U73 ( .A(FORWARDING__n417), .Y(FORWARDING__n264) );
  BUFx4f_ASAP7_75t_R FORWARDING___U74 ( .A(FORWARDING__n262), .Y(FORWARDING__n199) );
  BUFx3_ASAP7_75t_R FORWARDING___U75 ( .A(FORWARDING__n485), .Y(FORWARDING__n200) );
  HB1xp67_ASAP7_75t_R FORWARDING___U76 ( .A(FORWARDING__n201), .Y(FORWARDING__n177) );
  HB1xp67_ASAP7_75t_R FORWARDING___U77 ( .A(FORWARDING__n241), .Y(FORWARDING__n139) );
  HB1xp67_ASAP7_75t_R FORWARDING___U78 ( .A(FORWARDING__n140), .Y(FORWARDING__n241) );
  INVx1_ASAP7_75t_R FORWARDING___U79 ( .A(FORWARDING__n399), .Y(FORWARDING__n8) );
  AOI21xp5_ASAP7_75t_R FORWARDING___U80 ( .A1(FORWARDING__n17), .A2(FORWARDING__n18), .B(FORWARDING__n378), .Y(FORWARDING__n502) );
  INVx1_ASAP7_75t_R FORWARDING___U81 ( .A(FORWARDING__n242), .Y(FORWARDING__n18) );
  INVxp33_ASAP7_75t_R FORWARDING___U82 ( .A(FORWARDING__n184), .Y(forwarding_MEM_WB[12]) );
  AND2x2_ASAP7_75t_R FORWARDING___U83 ( .A(MEM_WB_mem_data[16]), .B(FORWARDING__n40), .Y(FORWARDING__FORWARDING__n407)
         );
  INVx2_ASAP7_75t_R FORWARDING___U84 ( .A(FORWARDING__n390), .Y(FORWARDING__n9) );
  AND2x4_ASAP7_75t_R FORWARDING___U85 ( .A(MEM_WB_mem_data[7]), .B(FORWARDING__n366), .Y(FORWARDING__n390)
         );
  INVxp33_ASAP7_75t_R FORWARDING___U86 ( .A(FORWARDING__n145), .Y(FORWARDING__n252) );
  HB1xp67_ASAP7_75t_R FORWARDING___U87 ( .A(FORWARDING__n477), .Y(FORWARDING__n145) );
  INVx1_ASAP7_75t_R FORWARDING___U88 ( .A(FORWARDING__n107), .Y(forwarding_MEM_WB[2]) );
  BUFx3_ASAP7_75t_R FORWARDING___U89 ( .A(FORWARDING__n436), .Y(FORWARDING__n193) );
  BUFx5_ASAP7_75t_R FORWARDING___U90 ( .A(FORWARDING__n368), .Y(FORWARDING__n372) );
  AND2x4_ASAP7_75t_R FORWARDING___U91 ( .A(MEM_WB_mem_data[15]), .B(FORWARDING__n368), .Y(FORWARDING__n405) );
  HB1xp67_ASAP7_75t_R FORWARDING___U92 ( .A(FORWARDING__n286), .Y(FORWARDING__n184) );
  BUFx2_ASAP7_75t_R FORWARDING___U93 ( .A(FORWARDING__n206), .Y(FORWARDING__n265) );
  HB1xp67_ASAP7_75t_R FORWARDING___U94 ( .A(FORWARDING__n495), .Y(FORWARDING__n206) );
  HB1xp67_ASAP7_75t_R FORWARDING___U95 ( .A(FORWARDING__n207), .Y(FORWARDING__n35) );
  HB1xp67_ASAP7_75t_R FORWARDING___U96 ( .A(FORWARDING__n185), .Y(FORWARDING__n286) );
  INVx2_ASAP7_75t_R FORWARDING___U97 ( .A(FORWARDING__n401), .Y(FORWARDING__n237) );
  HB1xp67_ASAP7_75t_R FORWARDING___U98 ( .A(FORWARDING__n360), .Y(FORWARDING__n371) );
  INVx4_ASAP7_75t_R FORWARDING___U99 ( .A(MEM_WB_mem_data[11]), .Y(FORWARDING__n21) );
  HB1xp67_ASAP7_75t_R FORWARDING___U100 ( .A(FORWARDING__n492), .Y(FORWARDING__n185) );
  HB1xp67_ASAP7_75t_R FORWARDING___U101 ( .A(FORWARDING__n2), .Y(forwarding_MEM_WB[30]) );
  AND2x2_ASAP7_75t_R FORWARDING___U102 ( .A(MEM_WB_mem_data[14]), .B(FORWARDING__n365), .Y(
        n403) );
  HB1xp67_ASAP7_75t_R FORWARDING___U103 ( .A(FORWARDING__n84), .Y(FORWARDING__n45) );
  INVx1_ASAP7_75t_R FORWARDING___U104 ( .A(FORWARDING__n376), .Y(FORWARDING__n10) );
  INVx3_ASAP7_75t_R FORWARDING___U105 ( .A(FORWARDING__n503), .Y(forwarding_MEM_WB[0]) );
  HB1xp67_ASAP7_75t_R FORWARDING___U106 ( .A(FORWARDING__n235), .Y(forwarding_MEM_WB[13]) );
  AO21x1_ASAP7_75t_R FORWARDING___U107 ( .A1(FORWARDING__n12), .A2(MEM_WB_ALU_result[10]), .B(
        n396), .Y(forwarding_MEM_WB[10]) );
  AND2x2_ASAP7_75t_R FORWARDING___U108 ( .A(MEM_WB_mem_data[10]), .B(FORWARDING__n365), .Y(
        n396) );
  BUFx12f_ASAP7_75t_R FORWARDING___U109 ( .A(FORWARDING__n373), .Y(FORWARDING__n57) );
  BUFx3_ASAP7_75t_R FORWARDING___U110 ( .A(FORWARDING__n491), .Y(FORWARDING__n70) );
  HB1xp67_ASAP7_75t_R FORWARDING___U111 ( .A(FORWARDING__n257), .Y(FORWARDING__n202) );
  INVxp33_ASAP7_75t_R FORWARDING___U112 ( .A(FORWARDING__n187), .Y(forwarding_MEM_WB[28]) );
  HB1xp67_ASAP7_75t_R FORWARDING___U113 ( .A(FORWARDING__n219), .Y(FORWARDING__n187) );
  HB1xp67_ASAP7_75t_R FORWARDING___U114 ( .A(FORWARDING__n500), .Y(FORWARDING__n257) );
  AND2x2_ASAP7_75t_R FORWARDING___U115 ( .A(MEM_WB_mem_data[4]), .B(FORWARDING__n369), .Y(FORWARDING__n384) );
  HB1xp67_ASAP7_75t_R FORWARDING___U116 ( .A(FORWARDING__n188), .Y(FORWARDING__n219) );
  INVx3_ASAP7_75t_R FORWARDING___U117 ( .A(FORWARDING__n487), .Y(forwarding_MEM_WB[17]) );
  HB1xp67_ASAP7_75t_R FORWARDING___U118 ( .A(FORWARDING__n252), .Y(forwarding_MEM_WB[29]) );
  BUFx3_ASAP7_75t_R FORWARDING___U119 ( .A(FORWARDING__n432), .Y(FORWARDING__n149) );
  HB1xp67_ASAP7_75t_R FORWARDING___U120 ( .A(FORWARDING__n478), .Y(FORWARDING__n188) );
  HB1xp67_ASAP7_75t_R FORWARDING___U121 ( .A(FORWARDING__n5), .Y(FORWARDING__n80) );
  INVx2_ASAP7_75t_R FORWARDING___U122 ( .A(FORWARDING__n148), .Y(FORWARDING__n254) );
  BUFx3_ASAP7_75t_R FORWARDING___U123 ( .A(FORWARDING__n409), .Y(FORWARDING__n285) );
  HB1xp67_ASAP7_75t_R FORWARDING___U124 ( .A(FORWARDING__n203), .Y(FORWARDING__n59) );
  AO21x1_ASAP7_75t_R FORWARDING___U125 ( .A1(FORWARDING__n23), .A2(FORWARDING__n24), .B(FORWARDING__n405), .Y(FORWARDING__n22) );
  NAND2xp5_ASAP7_75t_R FORWARDING___U126 ( .A(FORWARDING__n13), .B(FORWARDING__n14), .Y(FORWARDING__n15) );
  AND2x2_ASAP7_75t_R FORWARDING___U127 ( .A(FORWARDING__n15), .B(FORWARDING__n218), .Y(FORWARDING__n486) );
  INVx1_ASAP7_75t_R FORWARDING___U128 ( .A(FORWARDING__n217), .Y(FORWARDING__n13) );
  INVxp33_ASAP7_75t_R FORWARDING___U129 ( .A(FORWARDING__n360), .Y(FORWARDING__n14) );
  INVx1_ASAP7_75t_R FORWARDING___U130 ( .A(FORWARDING__n486), .Y(FORWARDING__n16) );
  INVxp33_ASAP7_75t_R FORWARDING___U131 ( .A(FORWARDING__n64), .Y(forwarding_MEM_WB[4]) );
  HB1xp67_ASAP7_75t_R FORWARDING___U132 ( .A(FORWARDING__n16), .Y(forwarding_MEM_WB[18]) );
  HB1xp67_ASAP7_75t_R FORWARDING___U133 ( .A(FORWARDING__n238), .Y(FORWARDING__n107) );
  HB1xp67_ASAP7_75t_R FORWARDING___U134 ( .A(FORWARDING__n247), .Y(FORWARDING__n198) );
  HB1xp67_ASAP7_75t_R FORWARDING___U135 ( .A(FORWARDING__n108), .Y(FORWARDING__n238) );
  HB1xp67_ASAP7_75t_R FORWARDING___U136 ( .A(FORWARDING__n501), .Y(FORWARDING__n108) );
  HB1xp67_ASAP7_75t_R FORWARDING___U137 ( .A(FORWARDING__n276), .Y(FORWARDING__n64) );
  HB1xp67_ASAP7_75t_R FORWARDING___U138 ( .A(FORWARDING__n194), .Y(FORWARDING__n110) );
  BUFx3_ASAP7_75t_R FORWARDING___U139 ( .A(FORWARDING__n57), .Y(FORWARDING__n367) );
  HB1xp67_ASAP7_75t_R FORWARDING___U140 ( .A(FORWARDING__n65), .Y(FORWARDING__n276) );
  BUFx3_ASAP7_75t_R FORWARDING___U141 ( .A(FORWARDING__n388), .Y(FORWARDING__n196) );
  HB1xp67_ASAP7_75t_R FORWARDING___U142 ( .A(FORWARDING__n111), .Y(FORWARDING__n194) );
  INVx1_ASAP7_75t_R FORWARDING___U143 ( .A(FORWARDING__n394), .Y(FORWARDING__n20) );
  BUFx2_ASAP7_75t_R FORWARDING___U144 ( .A(FORWARDING__n278), .Y(forwarding_MEM_WB[9]) );
  AND2x2_ASAP7_75t_R FORWARDING___U145 ( .A(FORWARDING__n234), .B(FORWARDING__n368), .Y(FORWARDING__n411) );
  HB1xp67_ASAP7_75t_R FORWARDING___U146 ( .A(FORWARDING__n141), .Y(FORWARDING__n140) );
  INVxp33_ASAP7_75t_R FORWARDING___U147 ( .A(FORWARDING__n240), .Y(FORWARDING__n109) );
  INVxp33_ASAP7_75t_R FORWARDING___U148 ( .A(FORWARDING__n136), .Y(forwarding_MEM_WB[5]) );
  BUFx3_ASAP7_75t_R FORWARDING___U149 ( .A(FORWARDING__n403), .Y(FORWARDING__n269) );
  HB1xp67_ASAP7_75t_R FORWARDING___U150 ( .A(FORWARDING__n112), .Y(FORWARDING__n111) );
  HB1xp67_ASAP7_75t_R FORWARDING___U151 ( .A(FORWARDING__n502), .Y(FORWARDING__n141) );
  HB1xp67_ASAP7_75t_R FORWARDING___U152 ( .A(FORWARDING__n66), .Y(FORWARDING__n65) );
  HB1xp67_ASAP7_75t_R FORWARDING___U153 ( .A(FORWARDING__n499), .Y(FORWARDING__n66) );
  HB1xp67_ASAP7_75t_R FORWARDING___U154 ( .A(FORWARDING__n497), .Y(FORWARDING__n112) );
  HB1xp67_ASAP7_75t_R FORWARDING___U155 ( .A(FORWARDING__n380), .Y(FORWARDING__n240) );
  INVxp33_ASAP7_75t_R FORWARDING___U156 ( .A(FORWARDING__n47), .Y(FORWARDING__n278) );
  HB1xp67_ASAP7_75t_R FORWARDING___U157 ( .A(FORWARDING__n299), .Y(FORWARDING__n224) );
  HB1xp67_ASAP7_75t_R FORWARDING___U158 ( .A(FORWARDING__n225), .Y(FORWARDING__n299) );
  HB1xp67_ASAP7_75t_R FORWARDING___U159 ( .A(FORWARDING__n204), .Y(FORWARDING__n33) );
  HB1xp67_ASAP7_75t_R FORWARDING___U160 ( .A(FORWARDING__n109), .Y(FORWARDING__n43) );
  HB1xp67_ASAP7_75t_R FORWARDING___U161 ( .A(FORWARDING__n494), .Y(FORWARDING__n47) );
  HB1xp67_ASAP7_75t_R FORWARDING___U162 ( .A(FORWARDING__n484), .Y(FORWARDING__n225) );
  HB1xp67_ASAP7_75t_R FORWARDING___U163 ( .A(FORWARDING__n226), .Y(FORWARDING__n179) );
  NOR2x1p5_ASAP7_75t_R FORWARDING___U164 ( .A(FORWARDING__n21), .B(FORWARDING__n23), .Y(FORWARDING__n397) );
  CKINVDCx20_ASAP7_75t_R FORWARDING___U165 ( .A(FORWARDING__FORWARDING__n244), .Y(FORWARDING__n24) );
  HB1xp67_ASAP7_75t_R FORWARDING___U166 ( .A(FORWARDING__n260), .Y(FORWARDING__n136) );
  INVxp33_ASAP7_75t_R FORWARDING___U167 ( .A(FORWARDING__n208), .Y(forwarding_MEM_WB[15]) );
  HB1xp67_ASAP7_75t_R FORWARDING___U168 ( .A(FORWARDING__n137), .Y(FORWARDING__n260) );
  INVxp33_ASAP7_75t_R FORWARDING___U169 ( .A(FORWARDING__n283), .Y(FORWARDING__n106) );
  HB1xp67_ASAP7_75t_R FORWARDING___U170 ( .A(FORWARDING__n429), .Y(FORWARDING__n283) );
  HB1xp67_ASAP7_75t_R FORWARDING___U171 ( .A(FORWARDING__n243), .Y(FORWARDING__n208) );
  BUFx3_ASAP7_75t_R FORWARDING___U172 ( .A(FORWARDING__n413), .Y(FORWARDING__n312) );
  HB1xp67_ASAP7_75t_R FORWARDING___U173 ( .A(FORWARDING__n138), .Y(FORWARDING__n137) );
  HB1xp67_ASAP7_75t_R FORWARDING___U174 ( .A(FORWARDING__n498), .Y(FORWARDING__n138) );
  BUFx3_ASAP7_75t_R FORWARDING___U175 ( .A(FORWARDING__n479), .Y(FORWARDING__n104) );
  HB1xp67_ASAP7_75t_R FORWARDING___U176 ( .A(FORWARDING__n489), .Y(FORWARDING__n243) );
  HB1xp67_ASAP7_75t_R FORWARDING___U177 ( .A(FORWARDING__n275), .Y(FORWARDING__n98) );
  HB1xp67_ASAP7_75t_R FORWARDING___U178 ( .A(FORWARDING__n106), .Y(FORWARDING__n26) );
  INVxp67_ASAP7_75t_R FORWARDING___U179 ( .A(FORWARDING__n142), .Y(forwarding_MEM_WB[7]) );
  HB1xp67_ASAP7_75t_R FORWARDING___U180 ( .A(FORWARDING__n231), .Y(FORWARDING__n142) );
  HB1xp67_ASAP7_75t_R FORWARDING___U181 ( .A(FORWARDING__n303), .Y(FORWARDING__n81) );
  BUFx3_ASAP7_75t_R FORWARDING___U182 ( .A(FORWARDING__n397), .Y(FORWARDING__n305) );
  HB1xp67_ASAP7_75t_R FORWARDING___U183 ( .A(FORWARDING__n144), .Y(FORWARDING__n143) );
  HB1xp67_ASAP7_75t_R FORWARDING___U184 ( .A(FORWARDING__n496), .Y(FORWARDING__n144) );
  HB1xp67_ASAP7_75t_R FORWARDING___U185 ( .A(FORWARDING__n143), .Y(FORWARDING__n231) );
  HB1xp67_ASAP7_75t_R FORWARDING___U186 ( .A(FORWARDING__n82), .Y(FORWARDING__n303) );
  HB1xp67_ASAP7_75t_R FORWARDING___U187 ( .A(FORWARDING__n493), .Y(FORWARDING__n82) );
  AND2x4_ASAP7_75t_R FORWARDING___U188 ( .A(MEM_WB_mem_data[20]), .B(FORWARDING__n367), .Y(
        n415) );
  HB1xp67_ASAP7_75t_R FORWARDING___U189 ( .A(FORWARDING__n83), .Y(FORWARDING__n28) );
  HB1xp67_ASAP7_75t_R FORWARDING___U190 ( .A(FORWARDING__n135), .Y(FORWARDING__n76) );
  BUFx3_ASAP7_75t_R FORWARDING___U191 ( .A(FORWARDING__n415), .Y(FORWARDING__n302) );
  HB1xp67_ASAP7_75t_R FORWARDING___U192 ( .A(FORWARDING__n10), .Y(FORWARDING__n181) );
  BUFx3_ASAP7_75t_R FORWARDING___U193 ( .A(FORWARDING__n104), .Y(FORWARDING__n281) );
  BUFx6f_ASAP7_75t_R FORWARDING___U194 ( .A(FORWARDING__n375), .Y(FORWARDING__n357) );
  BUFx2_ASAP7_75t_R FORWARDING___U195 ( .A(FORWARDING__n273), .Y(FORWARDING__n31) );
  BUFx3_ASAP7_75t_R FORWARDING___U196 ( .A(FORWARDING__n271), .Y(FORWARDING__n316) );
  INVx2_ASAP7_75t_R FORWARDING___U197 ( .A(FORWARDING__n490), .Y(forwarding_MEM_WB[14]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U198 ( .A(FORWARDING__n265), .Y(FORWARDING__n205) );
  INVx2_ASAP7_75t_R FORWARDING___U199 ( .A(FORWARDING__n205), .Y(forwarding_MEM_WB[8]) );
  BUFx6f_ASAP7_75t_R FORWARDING___U200 ( .A(FORWARDING__n85), .Y(FORWARDING__n61) );
  BUFx2_ASAP7_75t_R FORWARDING___U201 ( .A(FORWARDING__n279), .Y(FORWARDING__n49) );
  BUFx3_ASAP7_75t_R FORWARDING___U202 ( .A(FORWARDING__n51), .Y(FORWARDING__n50) );
  BUFx2_ASAP7_75t_R FORWARDING___U203 ( .A(FORWARDING__N29), .Y(FORWARDING__n51) );
  INVx1_ASAP7_75t_R FORWARDING___U204 ( .A(FORWARDING__n321), .Y(FORWARDING__n454) );
  BUFx2_ASAP7_75t_R FORWARDING___U205 ( .A(FORWARDING__n53), .Y(FORWARDING__n52) );
  BUFx2_ASAP7_75t_R FORWARDING___U206 ( .A(FORWARDING__n440), .Y(FORWARDING__n53) );
  BUFx4f_ASAP7_75t_R FORWARDING___U207 ( .A(FORWARDING__n438), .Y(FORWARDING__n54) );
  BUFx2_ASAP7_75t_R FORWARDING___U208 ( .A(FORWARDING__n462), .Y(FORWARDING__n55) );
  BUFx2_ASAP7_75t_R FORWARDING___U209 ( .A(FORWARDING__n444), .Y(FORWARDING__n56) );
  BUFx2_ASAP7_75t_R FORWARDING___U210 ( .A(FORWARDING__n87), .Y(FORWARDING__n60) );
  BUFx4f_ASAP7_75t_R FORWARDING___U211 ( .A(FORWARDING__n162), .Y(FORWARDING__n85) );
  BUFx3_ASAP7_75t_R FORWARDING___U212 ( .A(FORWARDING__n86), .Y(FORWARDING__n162) );
  BUFx2_ASAP7_75t_R FORWARDING___U213 ( .A(FORWARDING__N31), .Y(FORWARDING__n62) );
  BUFx2_ASAP7_75t_R FORWARDING___U214 ( .A(FORWARDING__n126), .Y(FORWARDING__n63) );
  INVx1_ASAP7_75t_R FORWARDING___U215 ( .A(FORWARDING__n384), .Y(FORWARDING__n67) );
  BUFx2_ASAP7_75t_R FORWARDING___U216 ( .A(FORWARDING__n456), .Y(FORWARDING__n68) );
  BUFx2_ASAP7_75t_R FORWARDING___U217 ( .A(FORWARDING__n507), .Y(FORWARDING__n69) );
  BUFx4f_ASAP7_75t_R FORWARDING___U218 ( .A(EX_MEM_ALU_result[24]), .Y(
        forwarding_EX_MEM[24]) );
  INVx1_ASAP7_75t_R FORWARDING___U219 ( .A(FORWARDING__n70), .Y(FORWARDING__n235) );
  BUFx3_ASAP7_75t_R FORWARDING___U220 ( .A(FORWARDING__n75), .Y(FORWARDING__n74) );
  BUFx2_ASAP7_75t_R FORWARDING___U221 ( .A(FORWARDING__n463), .Y(FORWARDING__n75) );
  BUFx4f_ASAP7_75t_R FORWARDING___U222 ( .A(FORWARDING__n74), .Y(FORWARDING__n223) );
  BUFx2_ASAP7_75t_R FORWARDING___U223 ( .A(FORWARDING__n113), .Y(FORWARDING__n78) );
  INVx1_ASAP7_75t_R FORWARDING___U224 ( .A(FORWARDING__n305), .Y(FORWARDING__n83) );
  INVx2_ASAP7_75t_R FORWARDING___U225 ( .A(FORWARDING__n398), .Y(FORWARDING__n304) );
  BUFx4f_ASAP7_75t_R FORWARDING___U226 ( .A(MEM_WB_ALU_result[11]), .Y(FORWARDING__n398) );
  INVx1_ASAP7_75t_R FORWARDING___U227 ( .A(FORWARDING__n193), .Y(FORWARDING__n84) );
  BUFx2_ASAP7_75t_R FORWARDING___U228 ( .A(FORWARDING__n481), .Y(FORWARDING__n86) );
  BUFx2_ASAP7_75t_R FORWARDING___U229 ( .A(FORWARDING__n460), .Y(FORWARDING__n88) );
  BUFx4f_ASAP7_75t_R FORWARDING___U230 ( .A(EX_MEM_ALU_result[16]), .Y(
        forwarding_EX_MEM[16]) );
  BUFx3_ASAP7_75t_R FORWARDING___U231 ( .A(FORWARDING__n90), .Y(FORWARDING__n89) );
  BUFx2_ASAP7_75t_R FORWARDING___U232 ( .A(FORWARDING__n443), .Y(FORWARDING__n90) );
  CKINVDCx10_ASAP7_75t_R FORWARDING___U233 ( .A(FORWARDING__n189), .Y(FORWARDING__n321) );
  BUFx4f_ASAP7_75t_R FORWARDING___U234 ( .A(EX_MEM_ALU_result[29]), .Y(
        forwarding_EX_MEM[29]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U235 ( .A(EX_MEM_ALU_result[23]), .Y(
        forwarding_EX_MEM[23]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U236 ( .A(EX_MEM_ALU_result[10]), .Y(
        forwarding_EX_MEM[10]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U237 ( .A(EX_MEM_ALU_result[2]), .Y(
        forwarding_EX_MEM[2]) );
  BUFx2_ASAP7_75t_R FORWARDING___U238 ( .A(FORWARDING__n449), .Y(FORWARDING__n92) );
  BUFx2_ASAP7_75t_R FORWARDING___U239 ( .A(FORWARDING__n446), .Y(FORWARDING__n93) );
  BUFx3_ASAP7_75t_R FORWARDING___U240 ( .A(FORWARDING__n95), .Y(FORWARDING__n94) );
  BUFx2_ASAP7_75t_R FORWARDING___U241 ( .A(FORWARDING__n459), .Y(FORWARDING__n95) );
  BUFx2_ASAP7_75t_R FORWARDING___U242 ( .A(FORWARDING__n450), .Y(FORWARDING__n102) );
  BUFx2_ASAP7_75t_R FORWARDING___U243 ( .A(FORWARDING__n282), .Y(FORWARDING__n105) );
  INVx1_ASAP7_75t_R FORWARDING___U244 ( .A(FORWARDING__n196), .Y(FORWARDING__n113) );
  BUFx2_ASAP7_75t_R FORWARDING___U245 ( .A(FORWARDING__n445), .Y(FORWARDING__n114) );
  BUFx2_ASAP7_75t_R FORWARDING___U246 ( .A(FORWARDING__n55), .Y(FORWARDING__n115) );
  BUFx3_ASAP7_75t_R FORWARDING___U247 ( .A(n62), .Y(FORWARDING__n229) );
  BUFx2_ASAP7_75t_R FORWARDING___U248 ( .A(FORWARDING__n488), .Y(FORWARDING__n116) );
  INVx1_ASAP7_75t_R FORWARDING___U249 ( .A(FORWARDING__n116), .Y(FORWARDING__n159) );
  BUFx6f_ASAP7_75t_R FORWARDING___U250 ( .A(FORWARDING__n119), .Y(FORWARDING__n118) );
  BUFx4f_ASAP7_75t_R FORWARDING___U251 ( .A(FORWARDING__n50), .Y(FORWARDING__n119) );
  OR2x2_ASAP7_75t_R FORWARDING___U252 ( .A(FORWARDING__n221), .B(FORWARDING__n454), .Y(FORWARDING__N29) );
  AND2x6_ASAP7_75t_R FORWARDING___U253 ( .A(FORWARDING__n120), .B(FORWARDING__n223), .Y(FORWARDING__n448) );
  BUFx2_ASAP7_75t_R FORWARDING___U254 ( .A(FORWARDING__n461), .Y(FORWARDING__n121) );
  BUFx4f_ASAP7_75t_R FORWARDING___U255 ( .A(EX_MEM_ALU_result[25]), .Y(
        forwarding_EX_MEM[25]) );
  BUFx2_ASAP7_75t_R FORWARDING___U256 ( .A(FORWARDING__N30), .Y(FORWARDING__n122) );
  BUFx2_ASAP7_75t_R FORWARDING___U257 ( .A(FORWARDING__n441), .Y(FORWARDING__n123) );
  BUFx2_ASAP7_75t_R FORWARDING___U258 ( .A(FORWARDING__n442), .Y(FORWARDING__n124) );
  OR3x1_ASAP7_75t_R FORWARDING___U259 ( .A(FORWARDING__n127), .B(FORWARDING__n114), .C(FORWARDING__n227), .Y(FORWARDING__n443) );
  INVx1_ASAP7_75t_R FORWARDING___U260 ( .A(FORWARDING__n89), .Y(FORWARDING__n125) );
  OR2x2_ASAP7_75t_R FORWARDING___U261 ( .A(FORWARDING__n54), .B(FORWARDING__n293), .Y(FORWARDING__N31) );
  INVx1_ASAP7_75t_R FORWARDING___U262 ( .A(FORWARDING__n62), .Y(FORWARDING__n126) );
  BUFx4f_ASAP7_75t_R FORWARDING___U263 ( .A(FORWARDING__n128), .Y(FORWARDING__n127) );
  BUFx3_ASAP7_75t_R FORWARDING___U264 ( .A(FORWARDING__n56), .Y(FORWARDING__n128) );
  BUFx4f_ASAP7_75t_R FORWARDING___U265 ( .A(EX_MEM_ALU_result[9]), .Y(
        forwarding_EX_MEM[9]) );
  BUFx2_ASAP7_75t_R FORWARDING___U266 ( .A(FORWARDING__N27), .Y(FORWARDING__n131) );
  BUFx2_ASAP7_75t_R FORWARDING___U267 ( .A(FORWARDING__n457), .Y(FORWARDING__n132) );
  BUFx2_ASAP7_75t_R FORWARDING___U268 ( .A(FORWARDING__n458), .Y(FORWARDING__n133) );
  OR3x1_ASAP7_75t_R FORWARDING___U269 ( .A(FORWARDING__n88), .B(FORWARDING__n248), .C(FORWARDING__n115), .Y(FORWARDING__n459) );
  INVx1_ASAP7_75t_R FORWARDING___U270 ( .A(FORWARDING__n94), .Y(FORWARDING__n134) );
  INVx1_ASAP7_75t_R FORWARDING___U271 ( .A(FORWARDING__n302), .Y(FORWARDING__n135) );
  BUFx4f_ASAP7_75t_R FORWARDING___U272 ( .A(EX_MEM_ALU_result[18]), .Y(
        forwarding_EX_MEM[18]) );
  BUFx2_ASAP7_75t_R FORWARDING___U273 ( .A(FORWARDING__n253), .Y(FORWARDING__n147) );
  BUFx3_ASAP7_75t_R FORWARDING___U274 ( .A(FORWARDING__n149), .Y(FORWARDING__n148) );
  BUFx2_ASAP7_75t_R FORWARDING___U275 ( .A(FORWARDING__n309), .Y(FORWARDING__n152) );
  BUFx3_ASAP7_75t_R FORWARDING___U276 ( .A(FORWARDING__n154), .Y(FORWARDING__n153) );
  BUFx2_ASAP7_75t_R FORWARDING___U277 ( .A(FORWARDING__n423), .Y(FORWARDING__n154) );
  BUFx4f_ASAP7_75t_R FORWARDING___U278 ( .A(EX_MEM_ALU_result[27]), .Y(
        forwarding_EX_MEM[27]) );
  BUFx3_ASAP7_75t_R FORWARDING___U279 ( .A(FORWARDING__n156), .Y(FORWARDING__n155) );
  BUFx2_ASAP7_75t_R FORWARDING___U280 ( .A(FORWARDING__n439), .Y(FORWARDING__n156) );
  BUFx3_ASAP7_75t_R FORWARDING___U281 ( .A(FORWARDING__n158), .Y(FORWARDING__n157) );
  BUFx2_ASAP7_75t_R FORWARDING___U282 ( .A(FORWARDING__n455), .Y(FORWARDING__n158) );
  BUFx4f_ASAP7_75t_R FORWARDING___U283 ( .A(n66), .Y(FORWARDING__n250) );
  OA21x2_ASAP7_75t_R FORWARDING___U284 ( .A1(FORWARDING__n160), .A2(FORWARDING__n360), .B(FORWARDING__n161), .Y(FORWARDING__n488) );
  BUFx4f_ASAP7_75t_R FORWARDING___U285 ( .A(MEM_WB_ALU_result[16]), .Y(FORWARDING__n408) );
  INVx2_ASAP7_75t_R FORWARDING___U286 ( .A(FORWARDING__n408), .Y(FORWARDING__n160) );
  INVx1_ASAP7_75t_R FORWARDING___U287 ( .A(FORWARDING__n407), .Y(FORWARDING__n161) );
  OA21x2_ASAP7_75t_R FORWARDING___U288 ( .A1(FORWARDING__n358), .A2(FORWARDING__n163), .B(FORWARDING__n60), .Y(FORWARDING__n481) );
  BUFx2_ASAP7_75t_R FORWARDING___U289 ( .A(FORWARDING__n426), .Y(FORWARDING__n163) );
  AND2x2_ASAP7_75t_R FORWARDING___U290 ( .A(MEM_WB_mem_data[25]), .B(FORWARDING__n374), .Y(
        n425) );
  BUFx2_ASAP7_75t_R FORWARDING___U291 ( .A(FORWARDING__N28), .Y(FORWARDING__n165) );
  BUFx2_ASAP7_75t_R FORWARDING___U292 ( .A(FORWARDING__n212), .Y(FORWARDING__n166) );
  BUFx4f_ASAP7_75t_R FORWARDING___U293 ( .A(n53), .Y(FORWARDING__n167) );
  BUFx4f_ASAP7_75t_R FORWARDING___U294 ( .A(n53), .Y(FORWARDING__n168) );
  BUFx2_ASAP7_75t_R FORWARDING___U295 ( .A(FORWARDING__n470), .Y(FORWARDING__n169) );
  BUFx4f_ASAP7_75t_R FORWARDING___U296 ( .A(n59), .Y(FORWARDING__n213) );
  BUFx4f_ASAP7_75t_R FORWARDING___U297 ( .A(n57), .Y(FORWARDING__n170) );
  BUFx4f_ASAP7_75t_R FORWARDING___U298 ( .A(n57), .Y(FORWARDING__n171) );
  BUFx4f_ASAP7_75t_R FORWARDING___U299 ( .A(FORWARDING__n464), .Y(FORWARDING__n172) );
  BUFx4f_ASAP7_75t_R FORWARDING___U300 ( .A(FORWARDING__n322), .Y(FORWARDING__n173) );
  BUFx4f_ASAP7_75t_R FORWARDING___U301 ( .A(FORWARDING__n323), .Y(FORWARDING__n174) );
  BUFx4f_ASAP7_75t_R FORWARDING___U302 ( .A(FORWARDING__n324), .Y(FORWARDING__n175) );
  AND2x6_ASAP7_75t_R FORWARDING___U303 ( .A(EX_MEM_RegWrite), .B(FORWARDING__n191), .Y(FORWARDING__n447) );
  INVx2_ASAP7_75t_R FORWARDING___U304 ( .A(FORWARDING__n172), .Y(FORWARDING__n191) );
  INVx4_ASAP7_75t_R FORWARDING___U305 ( .A(EX_MEM_rd[1]), .Y(FORWARDING__n469) );
  INVx2_ASAP7_75t_R FORWARDING___U306 ( .A(FORWARDING__n199), .Y(forwarding_MEM_WB[21]) );
  BUFx3_ASAP7_75t_R FORWARDING___U307 ( .A(FORWARDING__n200), .Y(FORWARDING__n262) );
  BUFx2_ASAP7_75t_R FORWARDING___U308 ( .A(FORWARDING__n472), .Y(FORWARDING__n183) );
  BUFx2_ASAP7_75t_R FORWARDING___U309 ( .A(FORWARDING__n287), .Y(FORWARDING__n186) );
  BUFx4f_ASAP7_75t_R FORWARDING___U310 ( .A(EX_MEM_ALU_result[20]), .Y(
        forwarding_EX_MEM[20]) );
  BUFx12f_ASAP7_75t_R FORWARDING___U311 ( .A(FORWARDING__n190), .Y(FORWARDING__n189) );
  BUFx12f_ASAP7_75t_R FORWARDING___U312 ( .A(FORWARDING__n447), .Y(FORWARDING__n190) );
  AND2x4_ASAP7_75t_R FORWARDING___U313 ( .A(FORWARDING__n174), .B(FORWARDING__n175), .Y(FORWARDING__n464) );
  AND2x4_ASAP7_75t_R FORWARDING___U314 ( .A(FORWARDING__n245), .B(FORWARDING__n466), .Y(FORWARDING__n322) );
  AND2x4_ASAP7_75t_R FORWARDING___U315 ( .A(FORWARDING__n307), .B(FORWARDING__n173), .Y(FORWARDING__n323) );
  AND2x4_ASAP7_75t_R FORWARDING___U316 ( .A(FORWARDING__n468), .B(FORWARDING__n469), .Y(FORWARDING__n324) );
  INVx6_ASAP7_75t_R FORWARDING___U317 ( .A(FORWARDING__n465), .Y(FORWARDING__n245) );
  OA21x2_ASAP7_75t_R FORWARDING___U318 ( .A1(FORWARDING__n360), .A2(FORWARDING__n192), .B(FORWARDING__n45), .Y(FORWARDING__n475) );
  BUFx2_ASAP7_75t_R FORWARDING___U319 ( .A(FORWARDING__n437), .Y(FORWARDING__n192) );
  AND2x2_ASAP7_75t_R FORWARDING___U320 ( .A(MEM_WB_mem_data[31]), .B(FORWARDING__n130), .Y(
        n436) );
  OA21x2_ASAP7_75t_R FORWARDING___U321 ( .A1(FORWARDING__n363), .A2(FORWARDING__n195), .B(FORWARDING__n78), .Y(FORWARDING__n497) );
  BUFx4f_ASAP7_75t_R FORWARDING___U322 ( .A(MEM_WB_ALU_result[6]), .Y(FORWARDING__n389) );
  INVx2_ASAP7_75t_R FORWARDING___U323 ( .A(FORWARDING__n389), .Y(FORWARDING__n195) );
  AND2x2_ASAP7_75t_R FORWARDING___U324 ( .A(MEM_WB_mem_data[6]), .B(FORWARDING__n369), .Y(FORWARDING__n388) );
  INVx1_ASAP7_75t_R FORWARDING___U325 ( .A(FORWARDING__n382), .Y(FORWARDING__n203) );
  INVx1_ASAP7_75t_R FORWARDING___U326 ( .A(FORWARDING__n269), .Y(FORWARDING__n204) );
  BUFx2_ASAP7_75t_R FORWARDING___U327 ( .A(FORWARDING__n392), .Y(FORWARDING__n267) );
  INVx1_ASAP7_75t_R FORWARDING___U328 ( .A(FORWARDING__n267), .Y(FORWARDING__n207) );
  BUFx2_ASAP7_75t_R FORWARDING___U329 ( .A(FORWARDING__n319), .Y(FORWARDING__n211) );
  OR2x2_ASAP7_75t_R FORWARDING___U330 ( .A(FORWARDING__n54), .B(FORWARDING__n288), .Y(FORWARDING__N28) );
  INVx1_ASAP7_75t_R FORWARDING___U331 ( .A(FORWARDING__n165), .Y(FORWARDING__n212) );
  BUFx3_ASAP7_75t_R FORWARDING___U332 ( .A(n59), .Y(FORWARDING__n214) );
  BUFx4f_ASAP7_75t_R FORWARDING___U333 ( .A(n60), .Y(FORWARDING__n215) );
  BUFx4f_ASAP7_75t_R FORWARDING___U334 ( .A(n60), .Y(FORWARDING__n216) );
  BUFx4f_ASAP7_75t_R FORWARDING___U335 ( .A(MEM_WB_ALU_result[18]), .Y(FORWARDING__n412) );
  INVx2_ASAP7_75t_R FORWARDING___U336 ( .A(FORWARDING__n412), .Y(FORWARDING__n217) );
  INVx1_ASAP7_75t_R FORWARDING___U337 ( .A(FORWARDING__n411), .Y(FORWARDING__n218) );
  OA21x2_ASAP7_75t_R FORWARDING___U338 ( .A1(FORWARDING__n357), .A2(FORWARDING__n220), .B(FORWARDING__n80), .Y(FORWARDING__n478) );
  BUFx2_ASAP7_75t_R FORWARDING___U339 ( .A(FORWARDING__n431), .Y(FORWARDING__n220) );
  BUFx12f_ASAP7_75t_R FORWARDING___U340 ( .A(FORWARDING__n222), .Y(FORWARDING__n221) );
  BUFx12f_ASAP7_75t_R FORWARDING___U341 ( .A(FORWARDING__n448), .Y(FORWARDING__n222) );
  AND2x4_ASAP7_75t_R FORWARDING___U342 ( .A(FORWARDING__n221), .B(FORWARDING__n321), .Y(FORWARDING__n438) );
  INVx1_ASAP7_75t_R FORWARDING___U343 ( .A(FORWARDING__n419), .Y(FORWARDING__n226) );
  BUFx4f_ASAP7_75t_R FORWARDING___U344 ( .A(FORWARDING__n228), .Y(FORWARDING__n227) );
  BUFx3_ASAP7_75t_R FORWARDING___U345 ( .A(FORWARDING__n93), .Y(FORWARDING__n228) );
  BUFx12f_ASAP7_75t_R FORWARDING___U346 ( .A(FORWARDING__n505), .Y(FORWARDING__n230) );
  OA21x2_ASAP7_75t_R FORWARDING___U347 ( .A1(FORWARDING__n361), .A2(FORWARDING__n232), .B(FORWARDING__n9), .Y(FORWARDING__n496) );
  BUFx2_ASAP7_75t_R FORWARDING___U348 ( .A(FORWARDING__n391), .Y(FORWARDING__n232) );
  BUFx2_ASAP7_75t_R FORWARDING___U349 ( .A(FORWARDING__n506), .Y(FORWARDING__n233) );
  BUFx6f_ASAP7_75t_R FORWARDING___U350 ( .A(MEM_WB_mem_data[18]), .Y(FORWARDING__n234) );
  OA21x2_ASAP7_75t_R FORWARDING___U351 ( .A1(FORWARDING__n236), .A2(FORWARDING__n359), .B(FORWARDING__n237), .Y(FORWARDING__n491) );
  BUFx2_ASAP7_75t_R FORWARDING___U352 ( .A(FORWARDING__n402), .Y(FORWARDING__n236) );
  OA21x2_ASAP7_75t_R FORWARDING___U353 ( .A1(FORWARDING__n364), .A2(FORWARDING__n239), .B(FORWARDING__n43), .Y(FORWARDING__n501) );
  BUFx2_ASAP7_75t_R FORWARDING___U354 ( .A(FORWARDING__n381), .Y(FORWARDING__n239) );
  AND2x2_ASAP7_75t_R FORWARDING___U355 ( .A(MEM_WB_mem_data[2]), .B(FORWARDING__n370), .Y(FORWARDING__n380) );
  BUFx2_ASAP7_75t_R FORWARDING___U356 ( .A(FORWARDING__n379), .Y(FORWARDING__n242) );
  BUFx12f_ASAP7_75t_R FORWARDING___U357 ( .A(EX_MEM_rd[3]), .Y(FORWARDING__n465) );
  BUFx2_ASAP7_75t_R FORWARDING___U358 ( .A(FORWARDING__n284), .Y(FORWARDING__n246) );
  INVx1_ASAP7_75t_R FORWARDING___U359 ( .A(FORWARDING__n285), .Y(FORWARDING__n247) );
  BUFx4f_ASAP7_75t_R FORWARDING___U360 ( .A(FORWARDING__n249), .Y(FORWARDING__n248) );
  BUFx3_ASAP7_75t_R FORWARDING___U361 ( .A(FORWARDING__n121), .Y(FORWARDING__n249) );
  BUFx3_ASAP7_75t_R FORWARDING___U362 ( .A(n66), .Y(FORWARDING__n251) );
  BUFx4f_ASAP7_75t_R FORWARDING___U363 ( .A(EX_MEM_ALU_result[6]), .Y(
        forwarding_EX_MEM[6]) );
  OA21x2_ASAP7_75t_R FORWARDING___U364 ( .A1(FORWARDING__n147), .A2(FORWARDING__n357), .B(FORWARDING__n254), .Y(FORWARDING__n477) );
  BUFx2_ASAP7_75t_R FORWARDING___U365 ( .A(MEM_WB_ALU_result[29]), .Y(FORWARDING__n433) );
  INVx1_ASAP7_75t_R FORWARDING___U366 ( .A(FORWARDING__n433), .Y(FORWARDING__n253) );
  BUFx4f_ASAP7_75t_R FORWARDING___U367 ( .A(FORWARDING__n256), .Y(ForwardB[0]) );
  BUFx3_ASAP7_75t_R FORWARDING___U368 ( .A(FORWARDING__n69), .Y(FORWARDING__n256) );
  OA21x2_ASAP7_75t_R FORWARDING___U369 ( .A1(FORWARDING__n363), .A2(FORWARDING__n258), .B(FORWARDING__n59), .Y(FORWARDING__n500) );
  BUFx2_ASAP7_75t_R FORWARDING___U370 ( .A(FORWARDING__n383), .Y(FORWARDING__n258) );
  AND2x2_ASAP7_75t_R FORWARDING___U371 ( .A(MEM_WB_mem_data[3]), .B(FORWARDING__n370), .Y(FORWARDING__n382) );
  OA21x2_ASAP7_75t_R FORWARDING___U372 ( .A1(FORWARDING__n364), .A2(FORWARDING__n259), .B(FORWARDING__n181), .Y(FORWARDING__n503) );
  BUFx2_ASAP7_75t_R FORWARDING___U373 ( .A(FORWARDING__n377), .Y(FORWARDING__n259) );
  AND2x2_ASAP7_75t_R FORWARDING___U374 ( .A(MEM_WB_mem_data[0]), .B(FORWARDING__n372), .Y(FORWARDING__n376) );
  OA21x2_ASAP7_75t_R FORWARDING___U375 ( .A1(FORWARDING__n363), .A2(FORWARDING__n261), .B(FORWARDING__n6), .Y(FORWARDING__n498) );
  BUFx4f_ASAP7_75t_R FORWARDING___U376 ( .A(MEM_WB_ALU_result[5]), .Y(FORWARDING__n387) );
  INVx2_ASAP7_75t_R FORWARDING___U377 ( .A(FORWARDING__n387), .Y(FORWARDING__n261) );
  OA21x2_ASAP7_75t_R FORWARDING___U378 ( .A1(FORWARDING__n97), .A2(FORWARDING__n263), .B(FORWARDING__n177), .Y(FORWARDING__n485) );
  BUFx4f_ASAP7_75t_R FORWARDING___U379 ( .A(MEM_WB_ALU_result[21]), .Y(FORWARDING__n418) );
  INVx2_ASAP7_75t_R FORWARDING___U380 ( .A(FORWARDING__n418), .Y(FORWARDING__n263) );
  AND2x2_ASAP7_75t_R FORWARDING___U381 ( .A(MEM_WB_mem_data[21]), .B(FORWARDING__n40), .Y(FORWARDING__n417) );
  OA21x2_ASAP7_75t_R FORWARDING___U382 ( .A1(FORWARDING__n362), .A2(FORWARDING__n266), .B(FORWARDING__n35), .Y(FORWARDING__n495) );
  BUFx2_ASAP7_75t_R FORWARDING___U383 ( .A(FORWARDING__n393), .Y(FORWARDING__n266) );
  AND2x2_ASAP7_75t_R FORWARDING___U384 ( .A(MEM_WB_mem_data[8]), .B(FORWARDING__n72), .Y(FORWARDING__n392)
         );
  OA21x2_ASAP7_75t_R FORWARDING___U385 ( .A1(FORWARDING__n359), .A2(FORWARDING__n268), .B(FORWARDING__n33), .Y(FORWARDING__n490) );
  BUFx2_ASAP7_75t_R FORWARDING___U386 ( .A(FORWARDING__n404), .Y(FORWARDING__n268) );
  BUFx2_ASAP7_75t_R FORWARDING___U387 ( .A(FORWARDING__n480), .Y(FORWARDING__n271) );
  BUFx2_ASAP7_75t_R FORWARDING___U388 ( .A(FORWARDING__n317), .Y(FORWARDING__n272) );
  INVx1_ASAP7_75t_R FORWARDING___U389 ( .A(FORWARDING__n427), .Y(FORWARDING__n273) );
  BUFx2_ASAP7_75t_R FORWARDING___U390 ( .A(FORWARDING__n311), .Y(FORWARDING__n274) );
  INVx1_ASAP7_75t_R FORWARDING___U391 ( .A(FORWARDING__n312), .Y(FORWARDING__n275) );
  BUFx4f_ASAP7_75t_R FORWARDING___U392 ( .A(EX_MEM_ALU_result[22]), .Y(
        forwarding_EX_MEM[22]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U393 ( .A(EX_MEM_ALU_result[15]), .Y(
        forwarding_EX_MEM[15]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U394 ( .A(EX_MEM_ALU_result[13]), .Y(
        forwarding_EX_MEM[13]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U395 ( .A(EX_MEM_ALU_result[7]), .Y(
        forwarding_EX_MEM[7]) );
  OA21x2_ASAP7_75t_R FORWARDING___U396 ( .A1(FORWARDING__n362), .A2(FORWARDING__n277), .B(FORWARDING__n67), .Y(FORWARDING__n499) );
  BUFx2_ASAP7_75t_R FORWARDING___U397 ( .A(FORWARDING__n385), .Y(FORWARDING__n277) );
  OA21x2_ASAP7_75t_R FORWARDING___U398 ( .A1(FORWARDING__n49), .A2(FORWARDING__n361), .B(FORWARDING__n20), .Y(FORWARDING__FORWARDING__n494) );
  BUFx2_ASAP7_75t_R FORWARDING___U399 ( .A(MEM_WB_ALU_result[9]), .Y(FORWARDING__n395) );
  INVx1_ASAP7_75t_R FORWARDING___U400 ( .A(FORWARDING__n395), .Y(FORWARDING__n279) );
  AND2x2_ASAP7_75t_R FORWARDING___U401 ( .A(MEM_WB_mem_data[9]), .B(FORWARDING__n366), .Y(FORWARDING__n394) );
  OA21x2_ASAP7_75t_R FORWARDING___U402 ( .A1(FORWARDING__FORWARDING__n357), .A2(FORWARDING__n280), .B(FORWARDING__n3), .Y(FORWARDING__n476) );
  BUFx2_ASAP7_75t_R FORWARDING___U403 ( .A(FORWARDING__n435), .Y(FORWARDING__n280) );
  OA21x2_ASAP7_75t_R FORWARDING___U404 ( .A1(FORWARDING__n105), .A2(FORWARDING__n358), .B(FORWARDING__n26), .Y(FORWARDING__n479) );
  BUFx2_ASAP7_75t_R FORWARDING___U405 ( .A(MEM_WB_ALU_result[27]), .Y(FORWARDING__n430) );
  INVx1_ASAP7_75t_R FORWARDING___U406 ( .A(FORWARDING__n430), .Y(FORWARDING__n282) );
  AND2x2_ASAP7_75t_R FORWARDING___U407 ( .A(MEM_WB_mem_data[27]), .B(FORWARDING__n371), .Y(
        n429) );
  OA21x2_ASAP7_75t_R FORWARDING___U408 ( .A1(FORWARDING__n246), .A2(FORWARDING__n360), .B(FORWARDING__n198), .Y(FORWARDING__n487) );
  BUFx2_ASAP7_75t_R FORWARDING___U409 ( .A(MEM_WB_ALU_result[17]), .Y(FORWARDING__n410) );
  INVx1_ASAP7_75t_R FORWARDING___U410 ( .A(FORWARDING__n410), .Y(FORWARDING__n284) );
  AND2x2_ASAP7_75t_R FORWARDING___U411 ( .A(MEM_WB_mem_data[17]), .B(FORWARDING__n366), .Y(
        n409) );
  OA21x2_ASAP7_75t_R FORWARDING___U412 ( .A1(FORWARDING__n186), .A2(FORWARDING__n358), .B(FORWARDING__n8), .Y(FORWARDING__n492) );
  BUFx2_ASAP7_75t_R FORWARDING___U413 ( .A(MEM_WB_ALU_result[12]), .Y(FORWARDING__n400) );
  INVx1_ASAP7_75t_R FORWARDING___U414 ( .A(FORWARDING__n400), .Y(FORWARDING__n287) );
  AND2x2_ASAP7_75t_R FORWARDING___U415 ( .A(MEM_WB_mem_data[12]), .B(FORWARDING__n129), .Y(
        n399) );
  BUFx6f_ASAP7_75t_R FORWARDING___U416 ( .A(FORWARDING__n289), .Y(FORWARDING__n288) );
  BUFx4f_ASAP7_75t_R FORWARDING___U417 ( .A(FORWARDING__n157), .Y(FORWARDING__n289) );
  BUFx2_ASAP7_75t_R FORWARDING___U418 ( .A(FORWARDING__n474), .Y(FORWARDING__n290) );
  BUFx2_ASAP7_75t_R FORWARDING___U419 ( .A(FORWARDING__n473), .Y(FORWARDING__n291) );
  BUFx2_ASAP7_75t_R FORWARDING___U420 ( .A(FORWARDING__n471), .Y(FORWARDING__n292) );
  BUFx6f_ASAP7_75t_R FORWARDING___U421 ( .A(FORWARDING__n294), .Y(FORWARDING__n293) );
  BUFx4f_ASAP7_75t_R FORWARDING___U422 ( .A(FORWARDING__n155), .Y(FORWARDING__n294) );
  BUFx2_ASAP7_75t_R FORWARDING___U423 ( .A(FORWARDING__n452), .Y(FORWARDING__n295) );
  BUFx2_ASAP7_75t_R FORWARDING___U424 ( .A(FORWARDING__n453), .Y(FORWARDING__n296) );
  BUFx2_ASAP7_75t_R FORWARDING___U425 ( .A(FORWARDING__n451), .Y(FORWARDING__n297) );
  BUFx6f_ASAP7_75t_R FORWARDING___U426 ( .A(n5), .Y(FORWARDING__n298) );
  OA21x2_ASAP7_75t_R FORWARDING___U427 ( .A1(FORWARDING__n359), .A2(FORWARDING__n300), .B(FORWARDING__n179), .Y(FORWARDING__n484) );
  BUFx2_ASAP7_75t_R FORWARDING___U428 ( .A(FORWARDING__n420), .Y(FORWARDING__n300) );
  AND2x2_ASAP7_75t_R FORWARDING___U429 ( .A(MEM_WB_mem_data[22]), .B(FORWARDING__n368), .Y(
        n419) );
  BUFx2_ASAP7_75t_R FORWARDING___U430 ( .A(FORWARDING__n416), .Y(FORWARDING__n301) );
  OA21x2_ASAP7_75t_R FORWARDING___U431 ( .A1(FORWARDING__n365), .A2(FORWARDING__n304), .B(FORWARDING__n28), .Y(FORWARDING__n493) );
  BUFx12f_ASAP7_75t_R FORWARDING___U432 ( .A(FORWARDING__n504), .Y(ForwardA[1]) );
  XNOR2x2_ASAP7_75t_R FORWARDING___U433 ( .A(ID_EX_rs1[4]), .B(FORWARDING__n466), .Y(FORWARDING__n471) );
  BUFx12f_ASAP7_75t_R FORWARDING___U434 ( .A(EX_MEM_rd[2]), .Y(FORWARDING__n467) );
  INVx5_ASAP7_75t_R FORWARDING___U435 ( .A(FORWARDING__n467), .Y(FORWARDING__n307) );
  BUFx4f_ASAP7_75t_R FORWARDING___U436 ( .A(EX_MEM_ALU_result[12]), .Y(
        forwarding_EX_MEM[12]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U437 ( .A(EX_MEM_ALU_result[8]), .Y(
        forwarding_EX_MEM[8]) );
  OA21x2_ASAP7_75t_R FORWARDING___U438 ( .A1(FORWARDING__n152), .A2(FORWARDING__n359), .B(FORWARDING__n310), .Y(FORWARDING__n482) );
  BUFx2_ASAP7_75t_R FORWARDING___U439 ( .A(MEM_WB_ALU_result[24]), .Y(FORWARDING__n424) );
  INVx1_ASAP7_75t_R FORWARDING___U440 ( .A(FORWARDING__n424), .Y(FORWARDING__n309) );
  AND2x2_ASAP7_75t_R FORWARDING___U441 ( .A(MEM_WB_mem_data[24]), .B(FORWARDING__n374), .Y(
        n423) );
  BUFx2_ASAP7_75t_R FORWARDING___U442 ( .A(MEM_WB_ALU_result[19]), .Y(FORWARDING__n414) );
  INVx1_ASAP7_75t_R FORWARDING___U443 ( .A(FORWARDING__n414), .Y(FORWARDING__n311) );
  AND2x2_ASAP7_75t_R FORWARDING___U444 ( .A(n24), .B(FORWARDING__n368), .Y(
        n413) );
  XOR2x2_ASAP7_75t_R FORWARDING___U445 ( .A(n52), .B(FORWARDING__n215), .Y(FORWARDING__n445) );
  XOR2x2_ASAP7_75t_R FORWARDING___U446 ( .A(n33), .B(FORWARDING__n167), .Y(FORWARDING__n446) );
  XNOR2x2_ASAP7_75t_R FORWARDING___U447 ( .A(FORWARDING__n213), .B(FORWARDING__n307), .Y(FORWARDING__n470) );
  XOR2x2_ASAP7_75t_R FORWARDING___U448 ( .A(n52), .B(FORWARDING__n214), .Y(FORWARDING__n461) );
  BUFx12f_ASAP7_75t_R FORWARDING___U449 ( .A(FORWARDING__n230), .Y(ForwardA[0]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U450 ( .A(EX_MEM_ALU_result[21]), .Y(
        forwarding_EX_MEM[21]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U451 ( .A(EX_MEM_ALU_result[17]), .Y(
        forwarding_EX_MEM[17]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U452 ( .A(EX_MEM_ALU_result[5]), .Y(
        forwarding_EX_MEM[5]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U453 ( .A(FORWARDING__n315), .Y(ForwardB[1]) );
  BUFx3_ASAP7_75t_R FORWARDING___U454 ( .A(FORWARDING__n233), .Y(FORWARDING__n315) );
  OA21x2_ASAP7_75t_R FORWARDING___U455 ( .A1(FORWARDING__n272), .A2(FORWARDING__n358), .B(FORWARDING__n31), .Y(FORWARDING__n480) );
  BUFx2_ASAP7_75t_R FORWARDING___U456 ( .A(MEM_WB_ALU_result[26]), .Y(FORWARDING__n428) );
  INVx1_ASAP7_75t_R FORWARDING___U457 ( .A(FORWARDING__n428), .Y(FORWARDING__n317) );
  AND2x2_ASAP7_75t_R FORWARDING___U458 ( .A(MEM_WB_mem_data[26]), .B(FORWARDING__n370), .Y(
        n427) );
  OA21x2_ASAP7_75t_R FORWARDING___U459 ( .A1(FORWARDING__n211), .A2(FORWARDING__n359), .B(FORWARDING__n320), .Y(FORWARDING__n483) );
  BUFx2_ASAP7_75t_R FORWARDING___U460 ( .A(MEM_WB_ALU_result[23]), .Y(FORWARDING__n422) );
  INVx1_ASAP7_75t_R FORWARDING___U461 ( .A(FORWARDING__n422), .Y(FORWARDING__n319) );
  XNOR2x2_ASAP7_75t_R FORWARDING___U462 ( .A(FORWARDING__n250), .B(FORWARDING__n468), .Y(FORWARDING__n473) );
  XNOR2x2_ASAP7_75t_R FORWARDING___U463 ( .A(n62), .B(FORWARDING__n469), .Y(FORWARDING__n474) );
  XOR2x2_ASAP7_75t_R FORWARDING___U464 ( .A(n33), .B(FORWARDING__n229), .Y(FORWARDING__n462) );
  XNOR2x2_ASAP7_75t_R FORWARDING___U465 ( .A(ID_EX_rs2[3]), .B(n34), .Y(FORWARDING__n440) );
  XNOR2x2_ASAP7_75t_R FORWARDING___U466 ( .A(ID_EX_rs1[3]), .B(n34), .Y(FORWARDING__n456) );
  XNOR2x2_ASAP7_75t_R FORWARDING___U467 ( .A(ID_EX_rs1[3]), .B(FORWARDING__n245), .Y(FORWARDING__n472) );
  BUFx4f_ASAP7_75t_R FORWARDING___U468 ( .A(EX_MEM_ALU_result[31]), .Y(
        forwarding_EX_MEM[31]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U469 ( .A(EX_MEM_ALU_result[30]), .Y(
        forwarding_EX_MEM[30]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U470 ( .A(EX_MEM_ALU_result[28]), .Y(
        forwarding_EX_MEM[28]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U471 ( .A(EX_MEM_ALU_result[26]), .Y(
        forwarding_EX_MEM[26]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U472 ( .A(EX_MEM_ALU_result[19]), .Y(
        forwarding_EX_MEM[19]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U473 ( .A(EX_MEM_ALU_result[14]), .Y(
        forwarding_EX_MEM[14]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U474 ( .A(EX_MEM_ALU_result[11]), .Y(
        forwarding_EX_MEM[11]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U475 ( .A(EX_MEM_ALU_result[4]), .Y(
        forwarding_EX_MEM[4]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U476 ( .A(EX_MEM_ALU_result[3]), .Y(
        forwarding_EX_MEM[3]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U477 ( .A(EX_MEM_ALU_result[1]), .Y(
        forwarding_EX_MEM[1]) );
  BUFx4f_ASAP7_75t_R FORWARDING___U478 ( .A(EX_MEM_ALU_result[0]), .Y(
        forwarding_EX_MEM[0]) );
  XOR2x2_ASAP7_75t_R FORWARDING___U479 ( .A(ID_EX_rs2[4]), .B(EX_MEM_rd[4]), .Y(FORWARDING__n450) );
  XOR2x2_ASAP7_75t_R FORWARDING___U480 ( .A(ID_EX_rs2[3]), .B(EX_MEM_rd[3]), .Y(FORWARDING__n451) );
  XOR2x2_ASAP7_75t_R FORWARDING___U481 ( .A(FORWARDING__n216), .B(EX_MEM_rd[2]), .Y(FORWARDING__n449) );
  XOR2x2_ASAP7_75t_R FORWARDING___U482 ( .A(FORWARDING__n168), .B(EX_MEM_rd[1]), .Y(FORWARDING__n453) );
  XOR2x2_ASAP7_75t_R FORWARDING___U483 ( .A(FORWARDING__n171), .B(EX_MEM_rd[0]), .Y(FORWARDING__n452) );
  INVx4_ASAP7_75t_R FORWARDING___U484 ( .A(EX_MEM_rd[4]), .Y(FORWARDING__n466) );
  INVx4_ASAP7_75t_R FORWARDING___U485 ( .A(EX_MEM_rd[0]), .Y(FORWARDING__n468) );
  XOR2x2_ASAP7_75t_R FORWARDING___U486 ( .A(n12), .B(FORWARDING__n251), .Y(FORWARDING__n460) );
  XOR2x2_ASAP7_75t_R FORWARDING___U487 ( .A(n12), .B(FORWARDING__n170), .Y(FORWARDING__n444) );
  XNOR2x2_ASAP7_75t_R FORWARDING___U488 ( .A(ID_EX_rs1[4]), .B(n36), .Y(FORWARDING__n457) );
  XNOR2x2_ASAP7_75t_R FORWARDING___U489 ( .A(ID_EX_rs2[4]), .B(n36), .Y(FORWARDING__n441) );
  BUFx12f_ASAP7_75t_R FORWARDING___U490 ( .A(FORWARDING__n57), .Y(FORWARDING__n368) );
  INVx1_ASAP7_75t_R FORWARDING___U491 ( .A(MEM_WB_ALU_result[0]), .Y(FORWARDING__n377) );
  INVx1_ASAP7_75t_R FORWARDING___U492 ( .A(MEM_WB_ALU_result[2]), .Y(FORWARDING__n381) );
  INVx1_ASAP7_75t_R FORWARDING___U493 ( .A(MEM_WB_ALU_result[3]), .Y(FORWARDING__n383) );
  INVx1_ASAP7_75t_R FORWARDING___U494 ( .A(MEM_WB_ALU_result[4]), .Y(FORWARDING__n385) );
  INVx1_ASAP7_75t_R FORWARDING___U495 ( .A(MEM_WB_ALU_result[7]), .Y(FORWARDING__n391) );
  INVx1_ASAP7_75t_R FORWARDING___U496 ( .A(MEM_WB_ALU_result[8]), .Y(FORWARDING__n393) );
  INVx1_ASAP7_75t_R FORWARDING___U497 ( .A(MEM_WB_ALU_result[14]), .Y(FORWARDING__n404) );
  INVx1_ASAP7_75t_R FORWARDING___U498 ( .A(MEM_WB_ALU_result[20]), .Y(FORWARDING__n416) );
  INVx1_ASAP7_75t_R FORWARDING___U499 ( .A(MEM_WB_ALU_result[22]), .Y(FORWARDING__n420) );
  INVx1_ASAP7_75t_R FORWARDING___U500 ( .A(MEM_WB_ALU_result[25]), .Y(FORWARDING__n426) );
  INVx1_ASAP7_75t_R FORWARDING___U501 ( .A(MEM_WB_ALU_result[28]), .Y(FORWARDING__n431) );
  INVx1_ASAP7_75t_R FORWARDING___U502 ( .A(MEM_WB_ALU_result[30]), .Y(FORWARDING__n435) );
  INVx1_ASAP7_75t_R FORWARDING___U503 ( .A(MEM_WB_ALU_result[31]), .Y(FORWARDING__n437) );
  AND4x1_ASAP7_75t_R FORWARDING___U504 ( .A(FORWARDING__n52), .B(FORWARDING__n125), .C(FORWARDING__n124), .D(FORWARDING__n123), .Y(FORWARDING__N30) );
  OA21x2_ASAP7_75t_R FORWARDING___U505 ( .A1(FORWARDING__n321), .A2(FORWARDING__n293), .B(FORWARDING__n221), .Y(FORWARDING__n442) );
  OR5x1_ASAP7_75t_R FORWARDING___U506 ( .A(FORWARDING__n92), .B(FORWARDING__n102), .C(FORWARDING__n297), .D(FORWARDING__n295), .E(FORWARDING__n296), 
        .Y(FORWARDING__n439) );
  AND4x1_ASAP7_75t_R FORWARDING___U507 ( .A(FORWARDING__n68), .B(FORWARDING__n134), .C(FORWARDING__n133), .D(FORWARDING__n132), .Y(FORWARDING__N27) );
  OA21x2_ASAP7_75t_R FORWARDING___U508 ( .A1(FORWARDING__n288), .A2(FORWARDING__n321), .B(FORWARDING__n221), .Y(FORWARDING__n458) );
  OR5x1_ASAP7_75t_R FORWARDING___U509 ( .A(n34), .B(n36), .C(n52), .D(n12), .E(n33), .Y(FORWARDING__n463) );
  OR5x1_ASAP7_75t_R FORWARDING___U510 ( .A(FORWARDING__n169), .B(FORWARDING__n292), .C(FORWARDING__n183), .D(FORWARDING__n291), .E(FORWARDING__n290), 
        .Y(FORWARDING__n455) );

  NOR2x1p5_ASAP7_75t_R DATA_HAZARD___U1 ( .A(DATA_HAZARD__n13), .B(DATA_HAZARD__n10), .Y(stall) );
  NAND2xp33_ASAP7_75t_R DATA_HAZARD___U2 ( .A(DATA_HAZARD__n7), .B(DATA_HAZARD__n8), .Y(DATA_HAZARD__n21) );
  NAND2xp33_ASAP7_75t_R DATA_HAZARD___U3 ( .A(DATA_HAZARD__n6), .B(DATA_HAZARD__n5), .Y(DATA_HAZARD__n8) );
  NAND2xp5_ASAP7_75t_R DATA_HAZARD___U4 ( .A(DATA_HAZARD__n2), .B(DATA_HAZARD__n1), .Y(DATA_HAZARD__n4) );
  NAND2xp5_ASAP7_75t_R DATA_HAZARD___U5 ( .A(DATA_HAZARD__n3), .B(DATA_HAZARD__n4), .Y(DATA_HAZARD__n22) );
  INVx1_ASAP7_75t_R DATA_HAZARD___U6 ( .A(ID_EX_rd[2]), .Y(DATA_HAZARD__n2) );
  INVxp67_ASAP7_75t_R DATA_HAZARD___U7 ( .A(IF_ID_rs1[2]), .Y(DATA_HAZARD__n1) );
  XNOR2xp5_ASAP7_75t_R DATA_HAZARD___U8 ( .A(n40), .B(ID_EX_rd[2]), .Y(DATA_HAZARD__n17) );
  NAND2xp33_ASAP7_75t_R DATA_HAZARD___U9 ( .A(IF_ID_rs1[2]), .B(ID_EX_rd[2]), .Y(DATA_HAZARD__n3) );
  NAND2xp33_ASAP7_75t_R DATA_HAZARD___U10 ( .A(n45), .B(ID_EX_rd[0]), .Y(DATA_HAZARD__n7) );
  INVxp67_ASAP7_75t_R DATA_HAZARD___U11 ( .A(n45), .Y(DATA_HAZARD__n5) );
  INVxp33_ASAP7_75t_R DATA_HAZARD___U12 ( .A(ID_EX_rd[0]), .Y(DATA_HAZARD__n6) );
  XNOR2xp5_ASAP7_75t_R DATA_HAZARD___U13 ( .A(DATA_HAZARD__n15), .B(ID_EX_rd[3]), .Y(DATA_HAZARD__n19) );
  NAND5xp2_ASAP7_75t_R DATA_HAZARD___U14 ( .A(DATA_HAZARD__n18), .B(DATA_HAZARD__n15), .C(DATA_HAZARD__n17), .D(DATA_HAZARD__n16), .E(DATA_HAZARD__n19), .Y(
        n9) );
  AND2x2_ASAP7_75t_R DATA_HAZARD___U15 ( .A(DATA_HAZARD__n11), .B(DATA_HAZARD__n9), .Y(DATA_HAZARD__n10) );
  NAND5xp2_ASAP7_75t_R DATA_HAZARD___U16 ( .A(DATA_HAZARD__n24), .B(DATA_HAZARD__n23), .C(DATA_HAZARD__n21), .D(DATA_HAZARD__n20), .E(DATA_HAZARD__n22), .Y(
        n11) );
  XNOR2xp5_ASAP7_75t_R DATA_HAZARD___U17 ( .A(ID_EX_rd[4]), .B(n28), .Y(DATA_HAZARD__n18) );
  XNOR2xp5_ASAP7_75t_R DATA_HAZARD___U18 ( .A(ID_EX_rd[3]), .B(DATA_HAZARD__n25), .Y(DATA_HAZARD__n24) );
  XNOR2xp5_ASAP7_75t_R DATA_HAZARD___U19 ( .A(ID_EX_rd[1]), .B(n27), .Y(DATA_HAZARD__n15) );
  XNOR2xp5_ASAP7_75t_R DATA_HAZARD___U20 ( .A(n43), .B(ID_EX_rd[0]), .Y(DATA_HAZARD__n16) );
  XNOR2xp5_ASAP7_75t_R DATA_HAZARD___U21 ( .A(ID_EX_rd[4]), .B(n42), .Y(DATA_HAZARD__n23) );
  BUFx3_ASAP7_75t_R DATA_HAZARD___U22 ( .A(DATA_HAZARD__n14), .Y(DATA_HAZARD__n13) );
  XNOR2xp5_ASAP7_75t_R DATA_HAZARD___U23 ( .A(n30), .B(ID_EX_rd[1]), .Y(DATA_HAZARD__n20) );
  BUFx2_ASAP7_75t_R DATA_HAZARD___U24 ( .A(ID_EX_MemRead), .Y(DATA_HAZARD__n25) );
  INVx1_ASAP7_75t_R DATA_HAZARD___U25 ( .A(DATA_HAZARD__n25), .Y(DATA_HAZARD__n14) );
  BUFx3_ASAP7_75t_R U2 ( .A(IF_ID_rs1[3]), .Y(n25) );
  BUFx4f_ASAP7_75t_R U3 ( .A(IF_ID_rs1[4]), .Y(n42) );
  BUFx4f_ASAP7_75t_R U4 ( .A(IF_ID_rs2[0]), .Y(n108) );
  BUFx4f_ASAP7_75t_R U5 ( .A(IF_ID_rs2[1]), .Y(n38) );
  INVx1_ASAP7_75t_R U6 ( .A(n38), .Y(n41) );
  BUFx6f_ASAP7_75t_R U7 ( .A(WB_write_back_data[15]), .Y(n69) );
  BUFx2_ASAP7_75t_R U8 ( .A(WB_write_back_data[2]), .Y(n71) );
  HB1xp67_ASAP7_75t_R U9 ( .A(n51), .Y(n2) );
  INVx1_ASAP7_75t_R U10 ( .A(n112), .Y(n29) );
  INVxp67_ASAP7_75t_R U11 ( .A(WB_write_back_data[24]), .Y(n112) );
  BUFx3_ASAP7_75t_R U12 ( .A(WB_write_back_data[9]), .Y(n63) );
  HB1xp67_ASAP7_75t_R U13 ( .A(WB_write_back_data[22]), .Y(n72) );
  HB1xp67_ASAP7_75t_R U14 ( .A(n2), .Y(n3) );
  HB1xp67_ASAP7_75t_R U15 ( .A(MEM_WB_mem_data[13]), .Y(n5) );
  HB1xp67_ASAP7_75t_R U16 ( .A(MEM_WB_rd[3]), .Y(n4) );
  INVxp33_ASAP7_75t_R U17 ( .A(n27), .Y(n6) );
  INVxp67_ASAP7_75t_R U18 ( .A(n110), .Y(n109) );
  HB1xp67_ASAP7_75t_R U19 ( .A(IF_ID_inst[1]), .Y(n7) );
  BUFx2_ASAP7_75t_R U20 ( .A(WB_write_back_data[13]), .Y(n81) );
  BUFx3_ASAP7_75t_R U21 ( .A(ID_EX_inst_addr[14]), .Y(n58) );
  BUFx3_ASAP7_75t_R U22 ( .A(WB_write_back_data[28]), .Y(n48) );
  BUFx2_ASAP7_75t_R U23 ( .A(ID_EX_inst_addr[7]), .Y(n56) );
  BUFx2_ASAP7_75t_R U24 ( .A(WB_write_back_data[29]), .Y(n64) );
  HB1xp67_ASAP7_75t_R U25 ( .A(MEM_WB_rd[0]), .Y(n8) );
  INVx1_ASAP7_75t_R U26 ( .A(n17), .Y(n18) );
  BUFx6f_ASAP7_75t_R U27 ( .A(WB_write_back_data[19]), .Y(n111) );
  BUFx2_ASAP7_75t_R U28 ( .A(WB_write_back_data[1]), .Y(n70) );
  BUFx3_ASAP7_75t_R U29 ( .A(WB_write_back_data[6]), .Y(n68) );
  HB1xp67_ASAP7_75t_R U30 ( .A(n42), .Y(n9) );
  BUFx4f_ASAP7_75t_R U31 ( .A(n21), .Y(n52) );
  INVxp67_ASAP7_75t_R U32 ( .A(WB_write_back_data[17]), .Y(n110) );
  INVx1_ASAP7_75t_R U33 ( .A(n41), .Y(n27) );
  BUFx3_ASAP7_75t_R U34 ( .A(WB_write_back_data[23]), .Y(n16) );
  HB1xp67_ASAP7_75t_R U35 ( .A(IF_ID_rs1[2]), .Y(n10) );
  BUFx3_ASAP7_75t_R U36 ( .A(MEM_WB_rd[2]), .Y(n51) );
  HB1xp67_ASAP7_75t_R U37 ( .A(WB_write_back_data[8]), .Y(n65) );
  BUFx2_ASAP7_75t_R U38 ( .A(WB_write_back_data[14]), .Y(n46) );
  INVxp33_ASAP7_75t_R U39 ( .A(n8), .Y(n11) );
  INVx1_ASAP7_75t_R U40 ( .A(n11), .Y(n12) );
  HB1xp67_ASAP7_75t_R U41 ( .A(IF_ID_rs2[2]), .Y(n40) );
  HB1xp67_ASAP7_75t_R U42 ( .A(MEM_WB_rd[4]), .Y(n13) );
  HB1xp67_ASAP7_75t_R U43 ( .A(MEM_WB_mem_data[25]), .Y(n14) );
  BUFx4f_ASAP7_75t_R U44 ( .A(IF_ID_rs2[3]), .Y(n31) );
  BUFx2_ASAP7_75t_R U45 ( .A(IF_ID_rs2[4]), .Y(n28) );
  HB1xp67_ASAP7_75t_R U46 ( .A(IF_ID_rs2[3]), .Y(n15) );
  BUFx3_ASAP7_75t_R U47 ( .A(WB_write_back_data[21]), .Y(n73) );
  INVxp33_ASAP7_75t_R U48 ( .A(n6), .Y(n44) );
  HB1xp67_ASAP7_75t_R U49 ( .A(ID_EX_inst_addr[16]), .Y(n39) );
  BUFx6f_ASAP7_75t_R U50 ( .A(WB_write_back_data[0]), .Y(n55) );
  INVx1_ASAP7_75t_R U51 ( .A(EX_read_reg_data_2[30]), .Y(n17) );
  INVx1_ASAP7_75t_R U52 ( .A(EX_read_reg_data_2[15]), .Y(n19) );
  INVxp67_ASAP7_75t_R U53 ( .A(n19), .Y(n20) );
  HB1xp67_ASAP7_75t_R U54 ( .A(IF_ID_rs1[1]), .Y(n30) );
  HB1xp67_ASAP7_75t_R U55 ( .A(n3), .Y(n21) );
  BUFx6f_ASAP7_75t_R U56 ( .A(WB_write_back_data[26]), .Y(n49) );
  BUFx6f_ASAP7_75t_R U57 ( .A(ID_EX_inst_addr[15]), .Y(n67) );
  INVxp67_ASAP7_75t_R U58 ( .A(EX_branch_addr[25]), .Y(n22) );
  INVxp67_ASAP7_75t_R U59 ( .A(n22), .Y(n23) );
  BUFx3_ASAP7_75t_R U60 ( .A(WB_write_back_data[7]), .Y(n61) );
  HB1xp67_ASAP7_75t_R U61 ( .A(MEM_WB_mem_data[19]), .Y(n24) );
  HB1xp67_ASAP7_75t_R U62 ( .A(n28), .Y(n26) );
  BUFx12f_ASAP7_75t_R U63 ( .A(n48), .Y(n47) );
  INVxp33_ASAP7_75t_R U64 ( .A(MEM_WB_rd[1]), .Y(n32) );
  INVx1_ASAP7_75t_R U65 ( .A(n32), .Y(n33) );
  HB1xp67_ASAP7_75t_R U66 ( .A(IF_ID_rs1[0]), .Y(n45) );
  HB1xp67_ASAP7_75t_R U67 ( .A(n4), .Y(n34) );
  INVx2_ASAP7_75t_R U68 ( .A(n37), .Y(n35) );
  INVx4_ASAP7_75t_R U69 ( .A(n35), .Y(n36) );
  BUFx4f_ASAP7_75t_R U70 ( .A(n54), .Y(n37) );
  HB1xp67_ASAP7_75t_R U71 ( .A(IF_ID_rs2[0]), .Y(n43) );
  HB1xp67_ASAP7_75t_R U72 ( .A(n13), .Y(n54) );
  BUFx12f_ASAP7_75t_R U73 ( .A(ID_EX_inst_14_), .Y(n50) );
  BUFx6f_ASAP7_75t_R U74 ( .A(ID_EX_rs2[1]), .Y(n53) );
  BUFx6f_ASAP7_75t_R U75 ( .A(ID_EX_rs2[0]), .Y(n57) );
  BUFx6f_ASAP7_75t_R U76 ( .A(ID_EX_rs1[2]), .Y(n59) );
  BUFx6f_ASAP7_75t_R U77 ( .A(ID_EX_rs2[2]), .Y(n60) );
  BUFx6f_ASAP7_75t_R U78 ( .A(ID_EX_rs1[1]), .Y(n62) );
  BUFx6f_ASAP7_75t_R U79 ( .A(ID_EX_rs1[0]), .Y(n66) );
  HB1xp67_ASAP7_75t_R U80 ( .A(EX_MEM_read_reg_data_2[30]), .Y(n74) );
  HB1xp67_ASAP7_75t_R U81 ( .A(EX_MEM_read_reg_data_2[28]), .Y(n75) );
  HB1xp67_ASAP7_75t_R U82 ( .A(EX_MEM_read_reg_data_2[19]), .Y(n76) );
  HB1xp67_ASAP7_75t_R U83 ( .A(EX_MEM_read_reg_data_2[14]), .Y(n77) );
  HB1xp67_ASAP7_75t_R U84 ( .A(EX_MEM_read_reg_data_2[11]), .Y(n78) );
  HB1xp67_ASAP7_75t_R U85 ( .A(EX_MEM_read_reg_data_2[3]), .Y(n79) );
  HB1xp67_ASAP7_75t_R U86 ( .A(EX_MEM_read_reg_data_2[1]), .Y(n80) );
  HB1xp67_ASAP7_75t_R U87 ( .A(EX_MEM_read_reg_data_2[15]), .Y(n82) );
  HB1xp67_ASAP7_75t_R U88 ( .A(EX_MEM_read_reg_data_2[13]), .Y(n83) );
  HB1xp67_ASAP7_75t_R U89 ( .A(EX_MEM_read_reg_data_2[12]), .Y(n84) );
  HB1xp67_ASAP7_75t_R U90 ( .A(EX_MEM_read_reg_data_2[10]), .Y(n85) );
  HB1xp67_ASAP7_75t_R U91 ( .A(EX_MEM_read_reg_data_2[9]), .Y(n86) );
  HB1xp67_ASAP7_75t_R U92 ( .A(EX_MEM_read_reg_data_2[8]), .Y(n87) );
  HB1xp67_ASAP7_75t_R U93 ( .A(EX_MEM_read_reg_data_2[7]), .Y(n88) );
  HB1xp67_ASAP7_75t_R U94 ( .A(EX_MEM_read_reg_data_2[6]), .Y(n89) );
  HB1xp67_ASAP7_75t_R U95 ( .A(EX_MEM_read_reg_data_2[5]), .Y(n90) );
  HB1xp67_ASAP7_75t_R U96 ( .A(EX_MEM_read_reg_data_2[4]), .Y(n91) );
  HB1xp67_ASAP7_75t_R U97 ( .A(EX_MEM_read_reg_data_2[2]), .Y(n92) );
  HB1xp67_ASAP7_75t_R U98 ( .A(EX_MEM_read_reg_data_2[0]), .Y(n93) );
  HB1xp67_ASAP7_75t_R U99 ( .A(EX_MEM_MemWrite), .Y(n94) );
  HB1xp67_ASAP7_75t_R U100 ( .A(EX_MEM_read_reg_data_2[31]), .Y(n95) );
  HB1xp67_ASAP7_75t_R U101 ( .A(EX_MEM_read_reg_data_2[29]), .Y(n96) );
  HB1xp67_ASAP7_75t_R U102 ( .A(EX_MEM_read_reg_data_2[27]), .Y(n97) );
  HB1xp67_ASAP7_75t_R U103 ( .A(EX_MEM_read_reg_data_2[26]), .Y(n98) );
  HB1xp67_ASAP7_75t_R U104 ( .A(EX_MEM_read_reg_data_2[25]), .Y(n99) );
  HB1xp67_ASAP7_75t_R U105 ( .A(EX_MEM_read_reg_data_2[24]), .Y(n100) );
  HB1xp67_ASAP7_75t_R U106 ( .A(EX_MEM_read_reg_data_2[23]), .Y(n101) );
  HB1xp67_ASAP7_75t_R U107 ( .A(EX_MEM_read_reg_data_2[22]), .Y(n102) );
  HB1xp67_ASAP7_75t_R U108 ( .A(EX_MEM_read_reg_data_2[21]), .Y(n103) );
  HB1xp67_ASAP7_75t_R U109 ( .A(EX_MEM_read_reg_data_2[20]), .Y(n104) );
  HB1xp67_ASAP7_75t_R U110 ( .A(EX_MEM_read_reg_data_2[18]), .Y(n105) );
  HB1xp67_ASAP7_75t_R U111 ( .A(EX_MEM_read_reg_data_2[17]), .Y(n106) );
  HB1xp67_ASAP7_75t_R U112 ( .A(EX_MEM_read_reg_data_2[16]), .Y(n107) );
endmodule
